(* synthesize *)
module sysInvalid_UInt_Dec ();
   Reg#(Bit#(4)) rg <- mkReg('d256);
endmodule
