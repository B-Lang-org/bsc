package CircPkg;

interface Ifc;
   method Bool m();
endinterface

endpackage
