package DataDefResGivenNum () where

data (Foo :: #) = Bar

