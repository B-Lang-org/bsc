module f(Action);
   (* foo *)
   action
      noAction;
   endaction
endmodule

