
(* prefix = "foo" *)
interface Ifc;
  method Bool start(Bool a, Bool b);
endinterface

