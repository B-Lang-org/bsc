import Methods::*;

(* noinline *)
function T add(T x, T y);
  return (x + y);
endfunction

