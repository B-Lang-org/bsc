function bit [3:0] f();
  bit [3:0] x;
  begin
    x = 3;
  end
  f = x;
endfunction
