(* synthesize *)
(* no_default_reset *)
module mkEUseDefaultReset();
   Reg#(Bit#(32)) r <- mkReg(0);
endmodule
