package RWire ;

// The entire contents of this package have been moved to the PreludeBSV package.

endpackage

