import ReExportTestDataConFull::*;

U#(Bool) u = Tag { b1: True, b2: False };
