package SizedLiteral where

x :: Bit 5
x = 5'd10
