typedef struct {
   t f;
} S#(type t);

