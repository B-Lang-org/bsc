import Vector::*;

(* synthesize *)
module sysRenameClock ( (* osc="O", gate="G" *)
                        Vector#(2,Clock) clks,
                        Empty ifc );
endmodule

