(* synthesize *)
module sysInvalid_Bit_Hex ();
   Reg#(Bit#(4)) rg <- mkReg('hFF);
endmodule
