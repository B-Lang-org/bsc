package ScopeInNestedWhens ( mkScopeInNestedWhens ) where

struct Foo =
    a :: Bit 5
    b :: Bit 6
  deriving (Bits)

mkScopeInNestedWhens :: Module Empty
mkScopeInNestedWhens =
    module
	r :: Reg (Bit 5)
	r <- mkRegU

	q :: Reg Foo
	q <- mkRegU

        rules
	    when (Foo { a; b }) <- q
	     rules {
	         when True
	           ==> r := zeroExtend a
	    }

	    when s <- r
	     rules {
	         when True
	           ==> r := s + 1
	    }
