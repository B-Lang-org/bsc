`define is 6
`define fs 6
`define full sysFromReal_6_6

`include "FromReal.bsv"
