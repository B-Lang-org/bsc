typedef union tagged {
   void First;
   void Second;
} TaggedUnionVoid;

