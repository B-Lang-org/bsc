module Banner();

initial
begin
  $display("Verilog testcase 1.0");
end

endmodule
