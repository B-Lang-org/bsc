package DegreePrimeVar1() where

a° :: a -> a
a° = id
