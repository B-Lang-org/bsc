typedef struct {
  int x;
  int y;
} Coord_t;

Coord_t coords;
coords.x = 1;
coords.y = 1;
