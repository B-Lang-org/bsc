
(* synthesize, doc="foo\nbar", doc="quux" *)
(* doc="glurph bloop" *)
module mkCommentOnModule ();
endmodule

