-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EBadExport2.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers an unbound export error (EBadExport)

-- Error Message : bsc EBadExport2.bs
-- bsc: Compilation errors:
-- "EBadExport2.bs", line 14, column 53, Unbound or multiply exported: "xyz"
-----------------------------------------------------------------------
package EBadExport2 (EBadExport2(..), mkEBadExport2, xyz) where

-- import Int

interface EBadExport2 =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32


mkEBadExport2 :: Module EBadExport2
mkEBadExport2 =
    module

        x :: Reg (Int 32)
        x <- mkReg 0

        y :: Reg (Int 32)
        y <- mkReg 0

        rules
          "Swap":
            when x > y, y /= 0
              ==> action
                      x := y
                      y := x

          "Subtract":
            when x <= y, y /= 0
              ==> action
                      y := y - x

        interface
            start ix iy = action
                              x := ix
                              y := iy
                          when y == 0
            result = x when y == 0
