module mkFoo();
  rule bogus;
    Bool x = True;
  endrule
endmodule

