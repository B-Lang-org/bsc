package DuplicateTypeParam_Interface_Classic where

interface Ifc a b a =
  m :: Action

