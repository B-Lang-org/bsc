import Prelude::*;