
interface Ifc;
  (* prefix="first", result="res", prefix="second" *)
  method Bool start(Bool a, Bool b);
endinterface

