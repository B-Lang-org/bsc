(* synthesize *)
module sysClockedBy_BadName (Clock c1,
			     (* clocked_by="foo" *) Bool b,
			     Clock c2,
			     Empty ifc);
endmodule

