
interface Ifc;
 (* result = "" *)
 method Bool check ();
endinterface

