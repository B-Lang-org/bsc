package Expr_Ap () where

x :: Bool
x = _ True False False

