(* synthesize *)
module sysDeriveResetClock_Unused #(Reset r2)();

endmodule
