(* reset_prefix="" *)
module sysEmptyRSTNAttrib ();
endmodule

