interface Ifc;
  method Action m();
  method Action m();
endinterface
