typedef union tagged {
   struct {
      Bool first;
      Bool second;
   } OneTwo;
   void Three;
} TaggedUnionStruct;
