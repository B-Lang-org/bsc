// Comment

`line(/file/path,4,foo,0)

Bool b = True;
