module sysRules2();
function Rules f();
   int fi=12;
   return fi;
endfunction

function Rules g();
   int gi=13;
   return gi;
endfunction
endmodule
