
(* synthesize *)
module mkTest();
   Reg#(Bit#(3)) rg <- mkReg(fromInteger(valueOf(8)));
endmodule
