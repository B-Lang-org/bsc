module test();
   Bool x = True;
   x[0] = False;
   Bool y = x;
endmodule

