
interface Ifc;
  (* port = "foo" *)
  method Action check (Bool x);
endinterface

