package Util;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

import Control::*;
import StmtFSM::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

interface Configs#(type a);
   interface Control cntrl;
   method a      _read();
endinterface

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

function String showBool (Bool value);
   if (value)
      return "True";
   else
      return "False";
endfunction

function a grab_left(b value)
   provisos(Bits#(a, sa), Bits#(b, sb), Add#(x, sa, sb));

   let zow = truncate(pack(value) >> fromInteger((valueOf(sb) - valueOf(sa))));

   return unpack(zow);
endfunction
   
function Integer getSizeOf(a value)
   provisos(Bits#(a, sa));
   return valueOf(sa);
endfunction

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

endpackage