export ǉiǉan;

// the lowercase lj digraph is neither uppercase nor titlecase, so ok for variable identifiers

function a ǉiǉan(a x);
    return id(x);
endfunction: ǉiǉan

