package CHasType () where

import List

x :: Bit a
x = fromInteger (length (Nil :: (List a)))
