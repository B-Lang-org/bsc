package TypeAliasParamGivenTooMany () where

type (Foo :: # -> # -> *) a = Bit a

