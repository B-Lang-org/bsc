
interface Ifc;
 (* ready = "ch eck" *)
 method Bool check ();
endinterface

