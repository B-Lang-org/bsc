package ReExportSame_TopGood;

import ReExportSame_Sub::*;

export ReExportSame_Sub::*;

endpackage
