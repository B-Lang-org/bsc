(* synthesize *)
module sysUndetRules();
   addRules(?);
endmodule

