function Bit#(1) f(Bit#(1) arr[], a idx);
   return (arr[idx]);
endfunction
