import Vector::*;

(* synthesize *)
module sysNameCollision ( Vector#(2,Bool) b,
                          Bool b_0,
                          Empty ifc);
endmodule

