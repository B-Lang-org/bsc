module mkFoo();
  Bool x;
  x = True;
endmodule

