import MultErrors1::*;

Module#(Empty) poisonTest = mkErrorTop;



