module sysCircularRegister(Empty);
  Reg#(Bool) r();
  mkReg#(r) the_r(r);
endmodule: sysCircularRegister

