typedef enum { Red, Blue, Green } Color;

Color c1 = Red;

Color c2 = Red(True,False);

