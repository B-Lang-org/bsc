function Action f();
  action
    bit[3:0] x;
    x = x;
  endaction
endfunction
