
function m#(t) fn()
provisos(Monad#(m));
  return (begin
          end);
endfunction
