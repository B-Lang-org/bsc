module sysAmbigTCon_SizeOf (Reg#(Bit#(SizeOf#(t))));
endmodule
