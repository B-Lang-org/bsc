`define size 4
`define modName sysTest4

`include "Test.bsv"

