package FromIntegerTooLarge ( ) where

sysFromIntegerTooLarge :: Module Empty
sysFromIntegerTooLarge =
    module
        reg :: Reg (Bit 1)
        reg <- mkReg 3
        rules
            when True
             ==> { reg := 3 }
