package DoubleClockPrefix where

{-# synthesize sysDoubleClockPrefix {
  gate_input_clocks = { default_clock },
  clock_prefix = "clk",
  clock_prefix = "c",
  gate_prefix = "gate",
  reset_prefix = "rst" } #-}
sysDoubleClockPrefix :: (IsModule m mType) => m Empty
sysDoubleClockPrefix = module
  r :: Reg (UInt 16) <- mkReg 0
  rules
    "test": when True ==>
      r := r + 1
