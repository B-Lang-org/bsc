Bit#(8) y = 0;

Bit#(8) x = truncate( zeroExtend (y) );

