Bit#(7) x = 72'b0000000;
