import Sub1::*;

(*synthesize*)
module mkTest (Ifc1);
endmodule

