package FieldSelectionFromDigit where

data T = T { bar :: Bool }

x :: Bool
x = 0.bar
