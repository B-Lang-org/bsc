typedef union tagged {
  struct {
     function a id(a in) id;
     Integer b;
  } MyId;
} Id;

