function Action f();
  action
    function bit[0:0] id(bit[0:0] x);
      return x;
    endfunction
  endaction
endfunction

