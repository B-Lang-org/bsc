`include `

