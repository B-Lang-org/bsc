(* synthesize *)
module sysUndet_SubModArg ();
  Reg#(Bit#(32)) rg <- mkReg(?);
endmodule
