function Action f();
  action
    bit[3:0] x;
    x = 5;
    x = x;
  endaction
endfunction
