-----------------------------------------------------------------------
-- Project: Bluespec

-- File: ENotAlwaysReady.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the ENotAlwaysReady error of the bluespec
-- compiler (Method not always ready {identifier})
--
-- Generates error when verilog code is requested for mkGCD
-----------------------------------------------------------------------


package ENotAlwaysReady () where

-- import Int

interface GCD =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32

{-# properties mkGCD = {
          alwaysReady
}#-}

mkGCD :: Module GCD
mkGCD =
    module
	x :: Reg (Int 32)
	x <- mkRegU

	y :: Reg (Int 32)
	y <- mkReg 0

        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0


