package VarDefn_Type () where

_ :: Bool
_ = True

