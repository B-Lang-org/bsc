package Expr_HasType () where

x :: Bool
x = (_ :: Bool)

