typedef Tuple2#(a,b)  T#(type a, type b, type a);
