package WFilePackageNameMismatch_Top() where

import WFilePackageNameMismatch_Sub
