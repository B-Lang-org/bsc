// These comments should not be lost

`define m(x) x

module sysTest();

`m(endmodule)

// more comments here
