module mkModIfc_TooManyArgs_TopLevel(Reg#(Bool,Bool));
endmodule
