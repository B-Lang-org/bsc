module mkFoo();
  Reg#(Bool) r;
  r <- mkRegU();
endmodule
