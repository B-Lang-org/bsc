(* noinline *)
function Maybe#(data_t) fnNoInline_Polymorphic(data_t x);
   return (Valid(x));
endfunction

