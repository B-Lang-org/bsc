import Vector::*;

(* synthesize *)
module sysVectorOutOfBounds1();
   Integer x[4] = {1, 2, 3, 4};
   Vector#(4, Integer) v = arrayToVector(x);
   Integer y = v[5];
   
   rule test;
      $display("%0d", y);
      $finish(0);
   endrule
   
endmodule
