module mkTest ();
  Bool b;
  Integer i;
  Bit#(8) v;
  {b,i,v} = tuple3(True,1,2);
endmodule
