export żuraw;
export gżegżółka;

function a żuraw(a x);
    return id(x);
endfunction: żuraw

function a gżegżółka(a x);
    return id(x);
endfunction: gżegżółka

