package StructComponentUse() where

import StructComponentDef
