package DupPkg;

Bool x = False;

endpackage
