package PackageEmptyNoTail;
endpackage
