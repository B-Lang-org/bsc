import Keywords::*;

Bool x = False;

