function bit[3:0] f();
  function bit[3:0] g(Bool x);
    g = 3;
  endfunction
  f = 3;
endfunction

