(* synthesize *)
module mkAbstractDeriveType();
   Type t = ?;
   messageM(printType(t));
endmodule
