package DataDefParamGivenNonNumUsedNum () where

data (Foo :: * -> *) a = Bar (Bit a)

