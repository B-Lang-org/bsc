function Action f();
  action
    Bool y;
    Bool x;
    x = y;
  endaction
endfunction
