(* synthesize *)
(* clock_prefix="always" *)
module sysCLKAttribVerilogKeyword ();
endmodule

