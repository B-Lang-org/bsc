package Expr () where

x :: Bool
x = _

