`define size 3
`define modName sysTest3

`include "Test.bsv"

