package WrongPkg;

Bool x = True;

endpackage

