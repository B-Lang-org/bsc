import DupPkg::*;

Bool z = x;

