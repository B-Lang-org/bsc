package NotDisplayable() where

data Test = A | B

foo :: Action
foo = $display A 