
`define m(x
