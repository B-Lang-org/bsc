import DeprecatedLibrary::*;

Bool x = myFunc(True);

