// Comment

`line(/file/path)

Bool b = True;

