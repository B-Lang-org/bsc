
(* descending_urgency = 1 *)
module sysT2();
endmodule

