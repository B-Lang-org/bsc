import "BVI" DisplayReal =
module vDisplayReal#(real r)(Empty ifc);
      
   port val = r;
   
endmodule
