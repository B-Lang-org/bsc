import DupObj::*;

Bool z = x;

