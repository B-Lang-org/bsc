// Valid attribute is wrong place

interface Foo ;
   method Action start () ;
      (* descending_urgency = 1 *)
   method Action stop () ;
endinterface

module sysT2();
endmodule

