
(* noinline=1, noinline=0 *)
function Bool testMultipleAttribFunc();
   return True;
endfunction

