import TestDataCon2::*;

function Bool myFn (U#(Bool) x1, U#(Bool) x2);
  return (x1 == x2);
endfunction

