module sysECtxIsModuleActionValue_AVBindInModBlock(Empty);
   let v <- $time;
   rule r;
      $display("World");
   endrule
endmodule
