typedef struct {
    Bit#(8) red;
    Bit#(16) red;
    Bit#(8) blue;
} RgbColor;
