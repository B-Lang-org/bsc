typeclass Extend#(type a, type b);
      function b grow(a x);
      function a shrink(b x);
endtypeclass: Extend