package Undet3(sysUndet3) where

sysUndet3 :: Module Empty
sysUndet3 =
  module
    x :: Reg (Bit 27) <- mkReg _
    counter :: Reg (Bit 16) <- mkReg 0

    rules
      when True ==> counter := counter + 1
      when True ==> if (counter < 16) then displayHex(x :: Bit 27) else $finish 0
