package EmptyAction_Braces where

a :: Action
a = action {}

x :: Integer
x = 17
