typedef enum { Red, Green, Blue } Color;

Color red;
red = Red;
