Real x = 1.57;
