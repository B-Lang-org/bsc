(* noinline *)
function Bit#(32) some_function(Bit#(32) foo);
   begin
      return(foo - 3);
   end
endfunction

