package DisjointRanges(sysDisjointRanges) where

import FIFO

-- Rules `foo' and `bar' conflict, as they both try to enq on q,
-- and are not logically disjoint.
-- The ADisjoint range checker erroneously concludes that they are.

sysDisjointRanges :: Module Empty
sysDisjointRanges =
    module
	a :: Reg (Bit 16) <- mkRegU
	b :: Reg Bool <- mkRegU
	c :: Reg Bool <- mkRegU
	d :: Reg (Bit 16) <- mkRegU
	q :: FIFO Bool <- mkFIFO
        rules
            "foo": when (a > 63 || b) && (not c && (d >= 10 && a <= 63))
	            ==> { q.enq True }
	    "bar": when True
	            ==> { q.enq False }
