bit [3:1] threeBits;
threeBits = 7;
