import TypeclassDupSuperAbstract_Wrapper::*;
import TypeclassDupSuperAbstract_Leaf::*;

function Bool fn(Bool x);
  return cmeth(x,True);
endfunction

