import Vector::*;
export Vector::*;
