module sysWrongLoc_InoutArg ((*osc="clk"*) Inout#(Bool) i, Empty e);
endmodule

