`define is 10
`define fs 10
`define full sysFromReal_10_10

`include "FromReal.bsv"
