import Vector::*;

(* synthesize *)
module sysNameCollision ( (* port="b" *)Vector#(2,Bool) xs,
                          Bool b_0,
                          Empty ifc);
endmodule

