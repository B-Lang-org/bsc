package Prefixes where

{-# synthesize sysPrefixes {
  gate_input_clocks = { default_clock },
  clock_prefix = "clk",
  gate_prefix = "gate",
  reset_prefix = "rst" } #-}
sysPrefixes :: (IsModule m mType) => m Empty
sysPrefixes = module
  r :: Reg (UInt 16) <- mkReg 0
  rules
    "test": when True ==>
      r := r + 1
