
interface Ifc;
 method Action check ((* port="arg" *)Bool x, (* port="arg" *)Bool y);
endinterface

