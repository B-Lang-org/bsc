package ETooGeneral where

x :: a
x = True

