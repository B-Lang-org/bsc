package Input;

typedef struct {Bit#(129) a;
                Bit#(129) b;
				Bit#(129) sum;
				Bit#(129) diff;
				Bit#(129) mult;
                Bit#(128) sum_127;
                Bit#(127) sum_126;
                Bit#(97) sum_96;
                Bit#(96) sum_95;
                Bit#(95) sum_94;
                Bit#(65) sum_64;
                Bit#(64) sum_63;
                Bit#(63) sum_62;
                Bit#(33) sum_32;
                Bit#(32) sum_31;
                Bit#(31) sum_30;
                Bit#(2) sum_1;
                Bit#(1) sum_0;
                Bit#(128) diff_127;
                Bit#(127) diff_126;
                Bit#(97) diff_96;
                Bit#(96) diff_95;
                Bit#(95) diff_94;
                Bit#(65) diff_64;
                Bit#(64) diff_63;
                Bit#(63) diff_62;
                Bit#(33) diff_32;
                Bit#(32) diff_31;
                Bit#(31) diff_30;
                Bit#(2) diff_1;
                Bit#(1) diff_0;
                Bit#(128) mult_127;
                Bit#(127) mult_126;
                Bit#(97) mult_96;
                Bit#(96) mult_95;
                Bit#(95) mult_94;
                Bit#(65) mult_64;
                Bit#(64) mult_63;
                Bit#(63) mult_62;
                Bit#(33) mult_32;
                Bit#(32) mult_31;
                Bit#(31) mult_30;
                Bit#(2) mult_1;
                Bit#(1) mult_0;
				Bit#(70) logical;} Inputs deriving(Bits,Eq);

endpackage : Input
