typedef struct { Bool f; } S;

