package StructComponentTop(sysStructComponentTop) where

import StructComponentUse

-- Compiling this should not cause an internal error.  The error
-- arises because StructComponentUse.bi includes instances for
-- SomeStruct°Cons2 but not the type declaration for it. (Bug #207).

sysStructComponentTop :: Module Empty
sysStructComponentTop = module {}
