import ExportAllExport::*;

Bool quux;
quux = foo || bar;
