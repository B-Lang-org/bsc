package SizedLiteralTest where

{-# verilog sysSizedLiteralTest #-}
sysSizedLiteralTest :: Module Empty
sysSizedLiteralTest =
  module
    let a :: Bit 17
        a = 17'h1_1_1
        b :: Bit 17
        b = 17'h111
        z :: Bit 17
	z = 273
        c :: UInt 4
	c = 4'b0__01_1_00
        d :: UInt 4
	d = 4'b001100
        y :: UInt 4
	y = 12
        e :: Int 12
	e = 12'o7_7_7_7
        f :: Int 12
	f = 12'o7777
        x :: Int 12
	x = (0 - 1)
    rules
      when True ==>
        action
	  $display "%b %b %b" (1'b0 ++ a) (2'b0 ++ b) (3'b0 ++ z)
          $display "%h %h %h" (4'b0 ++ pack c) (8'b0 ++ pack d) (12'b0 ++ pack y)
	  if a == b && b == z &&
	     c == d && d == y &&
	     e == f && f == x
	    then $display "PASS"
	    else $display "FAIL"
	  $finish 0
