(* synthesize *)
module sysOctalChars();
rule test;
$display("\000");
$display("\001");
$display("\002");
$display("\003");
$display("\004");
$display("\005");
$display("\006");
$display("\007");
$display("\010");
$display("\011");
$display("\012");
$display("\013");
$display("\014");
$display("\015");
$display("\016");
$display("\017");
$display("\020");
$display("\021");
$display("\022");
$display("\023");
$display("\024");
$display("\025");
$display("\026");
$display("\027");
$display("\030");
$display("\031");
$display("\032");
$display("\033");
$display("\034");
$display("\035");
$display("\036");
$display("\037");
$display("\040");
$display("\041");
$display("\042");
$display("\043");
$display("\044");
$display("\045");
$display("\046");
$display("\047");
$display("\050");
$display("\051");
$display("\052");
$display("\053");
$display("\054");
$display("\055");
$display("\056");
$display("\057");
$display("\060");
$display("\061");
$display("\062");
$display("\063");
$display("\064");
$display("\065");
$display("\066");
$display("\067");
$display("\070");
$display("\071");
$display("\072");
$display("\073");
$display("\074");
$display("\075");
$display("\076");
$display("\077");
$display("\100");
$display("\101");
$display("\102");
$display("\103");
$display("\104");
$display("\105");
$display("\106");
$display("\107");
$display("\110");
$display("\111");
$display("\112");
$display("\113");
$display("\114");
$display("\115");
$display("\116");
$display("\117");
$display("\120");
$display("\121");
$display("\122");
$display("\123");
$display("\124");
$display("\125");
$display("\126");
$display("\127");
$display("\130");
$display("\131");
$display("\132");
$display("\133");
$display("\134");
$display("\135");
$display("\136");
$display("\137");
$display("\140");
$display("\141");
$display("\142");
$display("\143");
$display("\144");
$display("\145");
$display("\146");
$display("\147");
$display("\150");
$display("\151");
$display("\152");
$display("\153");
$display("\154");
$display("\155");
$display("\156");
$display("\157");
$display("\160");
$display("\161");
$display("\162");
$display("\163");
$display("\164");
$display("\165");
$display("\166");
$display("\167");
$display("\170");
$display("\171");
$display("\172");
$display("\173");
$display("\174");
$display("\175");
$display("\176");
$display("\177");
$display("\200");
$display("\201");
$display("\202");
$display("\203");
$display("\204");
$display("\205");
$display("\206");
$display("\207");
$display("\210");
$display("\211");
$display("\212");
$display("\213");
$display("\214");
$display("\215");
$display("\216");
$display("\217");
$display("\220");
$display("\221");
$display("\222");
$display("\223");
$display("\224");
$display("\225");
$display("\226");
$display("\227");
$display("\230");
$display("\231");
$display("\232");
$display("\233");
$display("\234");
$display("\235");
$display("\236");
$display("\237");
$display("\240");
$display("\241");
$display("\242");
$display("\243");
$display("\244");
$display("\245");
$display("\246");
$display("\247");
$display("\250");
$display("\251");
$display("\252");
$display("\253");
$display("\254");
$display("\255");
$display("\256");
$display("\257");
$display("\260");
$display("\261");
$display("\262");
$display("\263");
$display("\264");
$display("\265");
$display("\266");
$display("\267");
$display("\270");
$display("\271");
$display("\272");
$display("\273");
$display("\274");
$display("\275");
$display("\276");
$display("\277");
$display("\300");
$display("\301");
$display("\302");
$display("\303");
$display("\304");
$display("\305");
$display("\306");
$display("\307");
$display("\310");
$display("\311");
$display("\312");
$display("\313");
$display("\314");
$display("\315");
$display("\316");
$display("\317");
$display("\320");
$display("\321");
$display("\322");
$display("\323");
$display("\324");
$display("\325");
$display("\326");
$display("\327");
$display("\330");
$display("\331");
$display("\332");
$display("\333");
$display("\334");
$display("\335");
$display("\336");
$display("\337");
$display("\340");
$display("\341");
$display("\342");
$display("\343");
$display("\344");
$display("\345");
$display("\346");
$display("\347");
$display("\350");
$display("\351");
$display("\352");
$display("\353");
$display("\354");
$display("\355");
$display("\356");
$display("\357");
$display("\360");
$display("\361");
$display("\362");
$display("\363");
$display("\364");
$display("\365");
$display("\366");
$display("\367");
$display("\370");
$display("\371");
$display("\372");
$display("\373");
$display("\374");
$display("\375");
$display("\376");
$display("\377");
endrule
endmodule
