import "BVI"
module mkMod(a);
   default_clock clk();
   default_reset rst();
endmodule

