import DupPkg::*;

Bool y = x;

