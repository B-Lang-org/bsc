package TypeAliasParamConflictingUses () where

data (Foo :: * -> *) a = Bar a

type Baz b = (Bit b, Foo b)

