import Vector::*;

module mkMod ();
   Reg#(Vector#(8,Integer)) rg <- mkRegU;
endmodule
