(* synthesize *)
module mkTest();
   Reg#(Bit#(TSub#(3,4))) rg <- mkRegU;
endmodule

