function Bool listy();
  Bool xsss[2][3][5];
  listy = xsss[0][2][4];
endfunction
