package CPrintType where

import List

class CPrintType a where
  cPrintType :: a -> String
  cPrintTypeP :: a -> String
  cPrintTypeP = cPrintType

instance (CPrintType a, CPrintTuple b) => CPrintType (a, b) where
  cPrintType _ = "(" +++ cPrintType (_ :: a) +++ ", " +++ cPrintTuple (_ :: b) +++ ")"

instance CPrintType () where
  cPrintType _ = "()"

class CPrintTuple a where
  cPrintTuple :: a -> String

instance (CPrintType a, CPrintTuple b) => CPrintTuple (a, b) where
  cPrintTuple _ = cPrintType (_ :: a) +++ ", " +++ cPrintTuple (_ :: b)

instance (CPrintType a) => CPrintTuple a where
  cPrintTuple = cPrintType

instance (Generic a r, CPrintType' r) => CPrintType a where
  cPrintType _ = cPrintType' (_ :: r)
  cPrintTypeP _ = cPrintTypeP' (_ :: r)

class CPrintType' a where
  cPrintType' :: a -> String
  cPrintTypeP' :: a -> String
  cPrintTypeP' = cPrintType'

instance CPrintType' (ConcPrim a) where
  cPrintType' _ = printType $ typeOf (_ :: a)

instance CPrintType' (Meta (MetaData n p () nc) r) where
  cPrintType' _ = stringOf n

instance (CPrintTypeArgs ta) => CPrintType' (Meta (MetaData n p ta nc) r) where
  cPrintType' _ = stringOf p +++ "." +++ stringOf n +++ " " +++ cPrintTypeArgs (_ :: ta)
  cPrintTypeP' _ = "(" +++ stringOf p +++ "." +++ stringOf n +++ " " +++ cPrintTypeArgs (_ :: ta) +++ ")"

class CPrintTypeArgs a where
  cPrintTypeArgs :: a -> String

instance (CPrintTypeArg a, CPrintTypeArgs b) => CPrintTypeArgs (a, b) where
  cPrintTypeArgs _ = cPrintTypeArg (_ :: a) +++ " " +++ cPrintTypeArgs (_ :: b)

instance (CPrintTypeArg a) => CPrintTypeArgs a where
  cPrintTypeArgs _ = cPrintTypeArg (_ :: a)

instance CPrintTypeArgs () where
  cPrintTypeArgs _ = ""

class CPrintTypeArg a where
  cPrintTypeArg :: a -> String

instance (CPrintType a) => CPrintTypeArg (StarArg a) where
  cPrintTypeArg _ = cPrintTypeP (_ :: a)

instance CPrintTypeArg (NumArg n) where
  cPrintTypeArg _ = integerToString $ valueOf n

instance CPrintTypeArg (StrArg s) where
  cPrintTypeArg _ = "\"" +++ stringOf s +++ "\""

instance (CPrintConType (c ())) => CPrintTypeArg (StarConArg c) where
  cPrintTypeArg _ = cPrintConType (_ :: c ())

instance (CPrintConType (c 0)) => CPrintTypeArg (NumConArg c) where
  cPrintTypeArg _ = cPrintConType (_ :: c 0)

instance CPrintTypeArg OtherConArg where
  cPrintTypeArg _ = "?"

class CPrintConType c where
  cPrintConType :: c -> String

instance (Generic c r, CPrintConType' r) => CPrintConType c where
  cPrintConType _ = cPrintConType' (_ :: r)

class CPrintConType' r where
  cPrintConType' :: r -> String

instance CPrintConType' (Meta (MetaData n p ta nc) r) where
  cPrintConType' _ = stringOf p +++ "." +++ stringOf n

instance (InitTuple (a, b) ta, CPrintTypeArgs ta) =>
    CPrintConType' (Meta (MetaData n p (a, b) nc) r) where
  cPrintConType' _ = "(" +++ stringOf p +++ "." +++ stringOf n +++
    " " +++ cPrintTypeArgs (_ :: ta) +++ ")"

class InitTuple a b | a -> b where {}
instance (InitTuple (b, c) d) => InitTuple (a, b, c) (a, d) where {}
instance InitTuple (a, b) a where {}

data Foo a b = A (UInt a)
             | B b Bool (Bit a)
             | C

data (Bar :: (* -> *) -> *) a = Bar (a Bool)
data (Baz :: (# -> *) -> (* -> * -> *) -> *) a b = Baz (a 42) (b Bool Integer)
data MyBit n = MyBit (Bit n)

sysCPrintType :: Module Empty
sysCPrintType = module
  rules
    when True ==> do
      $display (cPrintType (_ :: UInt 16))
      $display (cPrintType (_ :: (Either (Maybe Bool) String)))
      $display (cPrintType (_ :: (UInt 16, UInt 17)))
      $display (cPrintType (_ :: Foo 16 Real))
      $display (cPrintType $ from (_ :: Foo 16 Real))
      $display (cPrintType (_ :: Maybe (String, Integer)))
      $display (cPrintType (_ :: Bar Maybe))
      $display (cPrintType (_ :: Bar (Either Integer)))
      $display (cPrintType (_ :: Baz MyBit Either))
      $finish
