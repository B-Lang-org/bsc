package ResourceTwoRulesFail(sysResourceTwoRulesFail) where

import RegFile
import List

-- We are attempting to access six elements of an array simultaneously
-- in one rule, but Arrays only permit five simultaneous subs.
-- Expect to fail with a resource allocation error (unless
-- we compile with -resource-simple, in which case the compiler should
-- magically arbitrate between the two rules

type Index = Bit 8
type Value = Bit 8

lo :: Integer
lo = 0

hi :: Integer
hi = 2

lo2 :: Integer
lo2 = 10

hi2 :: Integer
hi2 = 12

sysResourceTwoRulesFail :: Module Empty
sysResourceTwoRulesFail =
      module
        r :: Reg Value
	r <- mkRegU
        s :: Reg Value
        s <- mkRegU
	a :: RegFile Index Value
	a <- mkRegFileFull
        rules
            "Bogus1":
               when True
                ==> r := (foldr (+) 0 $ map a.sub $ map fromInteger $ upto lo hi)
            "Bogus2":
               when True
                ==> s := (foldr (+) 0 $ map a.sub $ map fromInteger $ upto lo2 hi2)