function Bool listy();
  Bool xsss[2][3][5];
  listy = True;
endfunction
