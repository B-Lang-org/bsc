import TestDataConFull::*;

export U(..);

