module sysAmbigTCon_TMin (Reg#(Bit#(TMin#(x,y))));
endmodule
