
interface Ifc;
  interface Inout#(Bit#(32)) io_ifc;
endinterface

(*synthesize*)
module sysInoutProps_UnusedIfc (Ifc);
endmodule

