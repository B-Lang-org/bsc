
Bit#(0) x = 0'h0;

