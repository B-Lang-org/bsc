
module sysMultipleAttribRule();
   (* fire_when_enabled=1, fire_when_enabled=0 *)
   rule r;
      $display("Hi");
   endrule
endmodule

