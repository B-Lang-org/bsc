package ITransformConstantAcrossEquals ( ) where

sysITransformConstantAcrossEquals :: Module Empty
sysITransformConstantAcrossEquals =
    module
	r :: Reg (Bit 3) <- mkRegU
	x :: Reg (Bit 2) <- mkRegU
	y :: Reg (Bit 2) <- mkRegU
	z :: Reg (Bit 2) <- mkRegU

	rules
	  "Rule1":
	    when True ==>
	       action
		 if (r + 1 == 3) then x := x + 1 else x := x + 2
		 if (r - 1 == 3) then y := y + 1 else y := y + 2
		 if (((((r + 1) + 1) + 1) + 1) == 3)
		   then z := z + 1 else z := z + 2

	  "Rule2":
	    when True ==>
	       action
		 if (3 == r + 1) then x := x + 1 else x := x + 2
		 if (3 == r - 1) then y := y + 1 else y := y + 2
		 if (3 == ((((r + 1) + 1) + 1) + 1))
		   then z := z + 1 else z := z + 2

