import FieldDup_Wrapper::*;
import FieldDup_Leaf::*;

function Bool fn(S x);
  return x.f;
endfunction

