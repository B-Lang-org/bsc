package EmptyActionBreaks where

a :: Action
a = action

x :: Integer
x = 17
