typedef union tagged { Bool C; } U;
