module mkProvisoProvisoMismatch_Local();
   module mkMod(Reg#(t))
      provisos(Bits#(szt, j), Bits#(t, szt));
   endmodule
endmodule
