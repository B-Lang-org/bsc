function Bool fn(Bit#(n) x) provisos (Add#(2, k, n), Add#(n, k, 1));
   return ?;
endfunction

