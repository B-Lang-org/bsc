package Foreign () where

foreign _ :: Bit 1

