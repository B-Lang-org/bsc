////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

package ExtSDRAM;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

export mkExtSDRAM;

import RegFile::*;
import RegFile::*;
import SDRAM::*;

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

module mkExtSDRAM#(parameter ExtSDRAM ifc) (Empty);

   RegFile#(Bit#(AddrSize), Bit#(DataSize)) rom() ;
   mkRegFileLoad#("SRAM.handbuilt", 0, 'h1fffff) rom_inst(rom) ;

   rule every (True);
      action
	 if (ifc.rd && !ifc.wr)
	    begin
	       ifc.dOut( Valid(rom.sub(ifc.addr)) );
	    end
	 else 
	    ifc.dOut(Invalid);
      endaction
   endrule
   
endmodule

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

endpackage

////////////////////////////////////////////////////////////////////////////////
///
////////////////////////////////////////////////////////////////////////////////

