package ExportAllExport where

foo :: Bool
foo = True

bar :: Bool
bar = False
