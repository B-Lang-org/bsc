function Action f(Reg#(Bool) r);
  action
    r._write(True);
  endaction
endfunction

