function Bit#(1) f(Bit#(1) arr[], Bit#(a) idx);
  //provisos (PrimIndex#(Bit#(a)));
  //provisos (Add#(a,n,32));
   return (arr[idx]);
endfunction
