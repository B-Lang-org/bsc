package DataDefParamGivenNonNumUsedFunc () where

data (Foo :: * -> * -> *) x y = Bar (x y)

