import "BVI"
module mkFoo(i);
   Reg#(Bool) rg <- mkReg(True);
   // extra characters that cause the parser to stop parsing the module body
   );
   return ?;
endmodule
