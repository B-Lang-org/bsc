import List::*;

List#(Bool) xs = Prelude::Nil;
