
interface Ifc;
 (* enable = "always" *)
 method Action check ();
endinterface

(* synthesize *)
module mkKeyword (Ifc);
endmodule
