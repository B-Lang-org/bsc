package Math;

import Complex::*;
import FixedPoint::*;
import NumberTypes::*;
import Divide::*;
import SquareRoot::*;
import FloatingPoint::*;

// Re-export all imported packages
export Complex::*;
export FixedPoint::*;
export NumberTypes::*;
export Divide::*;
export SquareRoot::*;
export FloatingPoint::*;

endpackage
