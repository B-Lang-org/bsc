module mkFoo();
  Reg#(Bool) {x, y} ();
  mkReg#(True) the_r(x);
endmodule
