import Vector::*;

export Vector::*;
export replicateM;

