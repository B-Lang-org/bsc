module sysModDef_PortArg_Qmark(Bool ?, Empty ifc);
endmodule
