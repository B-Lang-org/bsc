interface Ifc;
  method Action m1(Bool s1, Bool s2);
endinterface

