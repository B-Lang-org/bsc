package Foo where

-- IMaybe creates separate ports for the valid bit and payload of a Maybe
-- at synthesis boundaries.
-- It deliberately does *not* derive Bits so that it isn't unexpectedly
-- packed or unpacked at synthesis boundaries.
interface IMaybe a =
    iValid :: Bool
    iValue :: a
  deriving(Eq)

iMaybe :: Maybe a -> IMaybe a
iMaybe ma = IMaybe { iValid = isValid ma; iValue = validValue ma }

data FooIn
  = Bar (Bit 2) (Maybe Bool)
  | Baz (UInt 5) (Int 7)
 deriving(Eq, Bits)

interface BarOut =
  bar_1 :: Bit 2
  bar_2 :: IMaybe Bool

interface BazOut =
  baz_1 :: UInt 5
  baz_2 :: Int 7

interface FooOut =
  bar :: IMaybe BarOut
  baz :: IMaybe BazOut

interface Foo =
  fooIn  :: FooIn -> Action {-# always_enabled #-}
  fooOut :: FooOut

{-# verilog mkFoo { noReady } #-}
mkFoo :: Module Foo
mkFoo = module
  fooWire <- mkBypassWire
  interface
    fooIn = fooWire._write
    fooOut = case fooWire of
               Bar bar_1 bar_2 ->
                  interface FooOut
                    bar = iMaybe $ Valid $ interface BarOut
                                             bar_1 = bar_1
                                             bar_2 = iMaybe bar_2
                    baz = iMaybe Invalid
               Baz baz_1 baz_2 ->
                  interface FooOut
                    bar = iMaybe Invalid
                    baz = iMaybe $ Valid $ interface BazOut
                                              baz_1 = baz_1
                                              baz_2 = baz_2