Bool _ = True;

// Test that "_" has type Bool by expecting a failure on mis-use
Bit#(8) y = _;

