import "BVI"
module mkMod(a#(Bit#(8)));
   default_clock clk();
   default_reset rst();
endmodule

