package TypeAliasPartialAppWithoutKindSig () where

type Foo = Bit

