(* synthesize, no_default_clock *)
module sysFixupRule_NoDefaultClock();
   rule r_disp;
      $display("Hello");
   endrule
endmodule
