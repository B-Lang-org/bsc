module mkProvisoBaseMismatch_TopLevel(Reg#(t))
   provisos(Add#(1,j,t));
endmodule
