// This should not compile because
// the parameter name is repeated
function Bool setInput(Bool x, Bool x);
    return False;
endfunction
