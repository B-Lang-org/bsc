package TypeAliasResGivenNonNumIsNum () where

type (Foo :: *) = 12

