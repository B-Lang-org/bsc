-- Tests to explore the compiler's output for derived Bits instances.
package DerivedBits where

interface TestTags =
  isA :: Bool
  isB :: Bool
  isC :: Bool
  isD :: Bool

data Orig = A (Bit 1)
          | B (Bit 1)
          | C (Bit 1)
          | D (Bit 1)
          deriving(Bits, Eq)

{-# verilog origReg #-}
origReg :: Module (Reg Orig)
origReg =
  module
    r <- mkRegU
    return r

{-# verilog origTest #-}
origTest :: Module TestTags
origTest =
  module
   r :: Reg Orig <- mkRegU
   interface TestTags
     isA = case r of
            A _ -> True
            _   -> False
     isB = case r of
            B _ -> True
            _   -> False
     isC = case r of
            C _ -> True
            _   -> False
     isD = case r of
            D _ -> True
            _   -> False

data Alt1 = A0
          | A1
          | B0
          | B1
          | C0
          | C1
          | D0
          | D1
  deriving(Bits)

{-# verilog altReg1 #-}
altReg1 :: Module (Reg Alt1)
altReg1 =
  module
    r <- mkRegU
    return r

{-# verilog alt1Test #-}
alt1Test :: Module TestTags
alt1Test =
  module
   r :: Reg Alt1 <- mkRegU
   interface TestTags
     isA = case r of
            A0  -> True
            A1  -> True
            _   -> False
     isB = case r of
            B0  -> True
            B1  -> True
            _   -> False
     isC = case r of
            C0  -> True
            C1  -> True
            _   -> False
     isD = case r of
            D0  -> True
            D1  -> True
            _   -> False

data Alt1a = A0
           | A1
           | B0
           | B1
           | C0
           | C1
  deriving(Bits)

{-# verilog altReg1a #-}
altReg1a :: Module (Reg Alt1a)
altReg1a =
  module
    r <- mkRegU
    return r

{-# verilog alt1aTest #-}
alt1aTest :: Module TestTags
alt1aTest =
  module
   r :: Reg Alt1 <- mkRegU
   interface TestTags
     isA = case r of
            A0  -> True
            A1  -> True
            _   -> False
     isB = case r of
            B0  -> True
            B1  -> True
            _   -> False
     isC = case r of
            C0  -> True
            C1  -> True
            _   -> False
     isD = False

data Alt2
    = A (Bit 1)
    | B (Bit 1)
    | C (Bit 1)
    | D
    deriving (Bits)

{-# verilog altReg2 #-}
altReg2 :: Module (Reg Alt2)
altReg2 =
  module
    r <- mkRegU
    return r

{-# verilog alt2Test #-}
alt2Test :: Module TestTags
alt2Test =
  module
   r :: Reg Alt2 <- mkRegU
   interface TestTags
     isA = case r of
            A _ -> True
            _   -> False
     isB = case r of
            B _ -> True
            _   -> False
     isC = case r of
            C _ -> True
            _   -> False
     isD = case r of
            D   -> True
            _   -> False

data Alt3
    = A (Bit 1)
    | B
    | C (Bit 1)
    | D (Bit 1)
    deriving (Bits)


{-# verilog altReg3 #-}
altReg3 :: Module (Reg Alt3)
altReg3 =
  module
    r <- mkRegU
    return r

{-# verilog alt3Test #-}
alt3Test :: Module TestTags
alt3Test =
  module
   r :: Reg Alt3 <- mkRegU
   interface TestTags
     isA = case r of
            A _ -> True
            _   -> False
     isB = case r of
            B   -> True
            _   -> False
     isC = case r of
            C _ -> True
            _   -> False
     isD = case r of
            D _ -> True
            _   -> False

data Tag4 = A | B | C | D
   deriving(Bits)

data Alt4 = Alt4 (Tag4, Bit 1)
  deriving(Bits)

{-# verilog altReg4 #-}
altReg4 :: Module (Reg Alt4)
altReg4 =
  module
    r <- mkRegU
    return r

{-# verilog alt4Test #-}
alt4Test :: Module TestTags
alt4Test =
  module
   r :: Reg Alt4 <- mkRegU
   interface TestTags
     isA = case r of
            Alt4 (A, _) -> True
            _           -> False
     isB = case r of
            Alt4 (B, _) -> True
            _           -> False
     isC = case r of
            Alt4 (C, _) -> True
            _           -> False
     isD = case r of
            Alt4 (D, _) -> True
            _           -> False

data Alt5
    = A (Bit 1)
    | B
    | C (Bit 1)
    | D
    deriving (Bits)

{-# verilog altReg5 #-}
altReg5 :: Module (Reg Alt5)
altReg5 =
  module
    r <- mkRegU
    return r

{-# verilog alt5Test #-}
alt5Test :: Module TestTags
alt5Test =
  module
   r :: Reg Alt5 <- mkRegU
   interface TestTags
     isA = case r of
            A _ -> True
            _   -> False
     isB = case r of
            B   -> True
            _   -> False
     isC = case r of
            C _ -> True
            _   -> False
     isD = case r of
            D   -> True
            _   -> False

data Alt6
    = A (Bit 1)
    | B (Bit 1)
    | C (Bit 1)
    deriving (Bits)

{-# verilog altReg6 #-}
altReg6 :: Module (Reg Alt6)
altReg6 =
  module
    r <- mkRegU
    return r

{-# verilog alt6Test #-}
alt6Test :: Module TestTags
alt6Test =
  module
   r :: Reg Alt6 <- mkRegU
   interface TestTags
     isA = case r of
            A _ -> True
            _   -> False
     isB = case r of
            B _ -> True
            _   -> False
     isC = case r of
            C _ -> True
            _   -> False
     isD = False

data C0 = E | F Orig | G C1
  deriving(Bits, Eq)

data C1 = H (UInt 2) (UInt 1) | I | J
  deriving(Bits, Eq)

interface TestTags2 =
  abcd :: TestTags
  isE :: Bool
  isF :: Bool
  isG :: Bool
  isH :: Bool
  isI :: Bool
  isJ :: Bool

{-# verilog c0Reg #-}
c0Reg :: Module (Reg C0)
c0Reg =
  module
    r <- mkRegU
    return r

{-# verilog c1Reg #-}
c1Reg :: Module (Reg C1)
c1Reg =
  module
    r <- mkRegU
    return r

{-# verilog c1Test #-}
c1Test :: Module TestTags2
c1Test =
  module
    r :: Reg C1 <- mkRegU
    interface
      abcd = interface TestTags
               isA = False
               isB = False
               isC = False
               isD = False
      isE = False
      isF = False
      isG = False
      isH = case r of
             H _ _ -> True
             _     -> False
      isI = r == I
      isJ = case r of
              J -> True
              _ -> False

{-# verilog c0Test #-}
c0Test :: Module TestTags2
c0Test =
  module
    r :: Reg C0 <- mkRegU
    interface
      abcd = interface TestTags
               isA = case r of
                       F (A _) -> True
                       _       -> False
               isB = case r of
                       F (B _) -> True
                       _       -> False
               isC = case r of
                       F (C _) -> True
                       _       -> False
               isD = case r of
                       F (D _) -> True
                       _       -> False
      isE = r == E
      isF = case r of
              F _ -> True
              _   -> False
      isG = case r of
              G _ -> True
              _   -> False
      isH = case r of
             G (H _ _) -> True
             _     -> False
      isI = r == (G I)
      isJ = case r of
              (G J) -> True
              _     -> False
