module mkTest1 (Empty);
    Reg#(Int#(32)) x();
    mkRegU#(1) the_x(x);
endmodule
