package ExportAllImport where

import ExportAllExport

quux :: Bool
quux = foo || bar
