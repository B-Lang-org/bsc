package Environment( ) where { }

