package StructDefParamGivenNonNumUsedNum () where

struct (Foo :: * -> *) a =
    bar :: Bit a

