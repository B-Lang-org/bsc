function Action f();
  action
    bit[3:0] x;
    x <- actionvalue return(3); endactionvalue;
  endaction
endfunction
