import List::*;

Prelude::List#(Prelude::Bool) xs = nil;
