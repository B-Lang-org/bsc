(* synthesize *)
module sysResetBy_BadName (Reset r1,
			   (* reset_by="foo" *) Bool b,
			   Reset r2,
			   Empty ifc);
endmodule

