module sysAmbigTCon_TMax (Reg#(Bit#(TMax#(x,y))));
endmodule
