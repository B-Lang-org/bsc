function Bool f() = False;
