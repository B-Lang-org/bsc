package Import1 (I) where
import Import0
interface I = m :: S
