import BasicReExport::*;
export BasicReExport::*;

