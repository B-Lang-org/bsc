(* synthesize *)
module sysInputPort#(Maybe#(Bool) test)(Empty);
endmodule
