package BindDummyDef () where

_ :: Int 32
_ = _

