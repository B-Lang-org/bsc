Rules rs;
rs = rules
       rule foo; endrule
       rule bar; endrule
     endrules;
