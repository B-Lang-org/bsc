package TypeAliasParamGivenTooFew_ToNone () where

type (Foo :: *) a = Bit a

