// Valid attribute is wrong place

interface Foo ;
   method Action start () ;
      (* result = "x1" *)
   interface Reg#(int)  rint ;
   method Action stop () ;
endinterface

module sysT2();
endmodule

