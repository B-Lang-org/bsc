
module BypassWire0();

endmodule
