export foo;

Bool foo;
foo = True;

Integer foo;
foo = 5;
