(* synthesize *)
(* gate_input_clocks = "default_clock" *)
module sysGateDefaultClock #(Clock c1, Clock c2, Clock c3) ();
endmodule

