(* synthesize *)
(* gate_all_clocks *)
module sysGateAllClocks #(Clock c1, Clock c2, Clock c3) ();
endmodule

