package SizedLiteralAmbig where

{-# verilog mkTop { no_default_reset } #-}
mkTop :: Module Empty
mkTop =
  module
    let a :: Bit 17
        a = 17'h1_1_1
        b = 17'h111
	z = 273
        c :: UInt 4
	c = 4'b0__01_1_00
	d = 4'b001100
	y = 12
        e :: Int 12
	e = 12'o7_7_7_7
	f = 12'o7777
	x = (0 - 1)
    rules
      when True ==>
        action
	  $display a " " c " " e
	  if a == b && b == z &&
	     c == d && d == y &&
	     e == f && f == x
	    then $display "PASS"
	    else $display "FAIL"
	  $finish 0
