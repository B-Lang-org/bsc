(* noinline *)
function Bool myAnd (Bool x, Bool y);
   return (x && y);
endfunction

