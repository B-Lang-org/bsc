package PackageModuleEmpty;
  module mkEmpty();
  endmodule: mkEmpty
endpackage: PackageModuleEmpty
