package TestExcludeOK where

import Exclude

d :: Integer
d = b + c
