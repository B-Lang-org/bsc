function Action f();
  Bool y;
  f = y;
endfunction
