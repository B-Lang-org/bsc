package DollarColonEqualsPrecedence1 where

foo :: Reg Bool -> Reg Bool
foo = id

bar :: Reg Bool -> Action
bar r = foo $ r := False

