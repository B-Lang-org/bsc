bit onebit;
onebit = 1;

bit [3:0] fourBits;
fourBits = 15;
