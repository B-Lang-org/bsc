
`undef - 

Bool x = True;

