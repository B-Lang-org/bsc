import DeprecatedLibrary::*;

Bool y = True;

