package Misc;

import Arbiter::*;
import BRAM::*;
import BRAMFIFO::*;
import BuildList::*;
import BuildVector::*;
import BUtils::*;
import BypassReg::*;
import Cntrs::*;
import DefaultValue ::*;
import Gray::*;
import GrayCounter::*;
import HList::*;
import Randomizable::*;
import SpecialFIFOs::*;
import AlignedFIFOs::*;
import TieOff ::*;
import DummyDriver ::*;
import Gearbox ::*;
import UnitAppendList::*;
import EdgeDetect::*;
import CRC::*;
import CommitIfc::*;
import NullCrossingFIFOF::*;
import MIMO::*;
import Memory::*;
import Arbitrate::*;
import Printf::*;
import PAClib::*;

endpackage
