function f(x, y);
  f = x || y;
endfunction: f
