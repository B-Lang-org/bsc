typeclass Foo#(type x)
 dependencies (x determines x);
   function Bool fooFn(x x1);
endtypeclass
