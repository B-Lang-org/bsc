package Contexts;

import ModuleContext::*;
import ModuleCollect::*;

// imported so that .bo files are generated
import CBus::*;
import LBus::*;



export ModuleContext::*;
export ModuleCollect::*;

endpackage
