----------------------------------------------------
-- FileName : MulticlockFIFO.bs
-- Author   : Interra
-- BugID    : 239
-- CommandLine : bsc -verilog -g mkTest MulticlockFIFO.bs
-- Status : Assigned
----------------------------------------------------

package MulticlockFIFO ( ) where

import ClockConv
import GetPut

mkMCFIFO :: (Bits a sa) => Clock -> Module (Closed (Get a), Put a)
mkMCFIFO clk2 =
     let mf :: Module (Closed (Get a), Put a)
         mf = module
                  (g, p) :: (Get a, Put a) <- mkGetPut
                  return (close g, p)

     in  clockConv clk2 mf

mkTest :: Clock -> Module (Closed (Get (Bit 5)), Put (Bit 5))
mkTest = mkMCFIFO
