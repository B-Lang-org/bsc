package TLMDefines;

typedef Bit#(8) TLMId;

endpackage
