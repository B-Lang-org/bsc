(* synthesize *)
(* no_default_clock *)
module mkEUseDefaultClock();
   Reg#(Bit#(32)) r <- mkRegU;
endmodule
