export とり;

// hiragana are not unicode uppercase letters

typedef union tagged {
   Bool つる
   void ふくろう;
} とり;

