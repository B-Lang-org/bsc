function Bool fn(Bool ?);
  return True;
endfunction
