
// User made a mistake in the syntax
`ifdef (verbosity >= 2)
Bool x = True;
`endif

