export foo;

Bool foo;
foo = True;
