typedef UInt#(8) Int;

function Int f(Int x, Int y);
   return x + y + 2;
endfunction

