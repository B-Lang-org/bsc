// This is quite contrived
typedef 4 ConstT#(numeric type a);

typedef Bit#(ConstT#(1)) Foo;

