import RightPkg::*;

Bool y = x;

