import List::*;

(* synthesize *)
module sysPrintType6();
   messageM(printType(typeOf(map)));
endmodule
