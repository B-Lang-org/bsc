package PackageEmpty;
endpackage: bogus
