package Defl_Clauses_NoType () where

x :: Bool
x = let _ 0 = True
        _ v = False
    in  True

