import Test:: *;

`include "IncDep1.bsv"
