function Action f(bit[3:0] x);
  action
    f(3);
  endaction
endfunction
