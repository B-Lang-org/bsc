package VarDefn_Clauses_NoType () where

_ 0 = True
_ v = False

