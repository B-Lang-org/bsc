-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EUnifyKind1.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers a Kind error (EUnifyKind)

-- Error Message : bsc EUnifyKind1.bs
-- bsc: Compilation errors:
-- "EUnifyKind1.bs", line 40, column 13, Kind error at:
-- Mystruct

-- Expected kind:
-- *

-- Inferred kind:
-- * -> *
-----------------------------------------------------------------------

package EUnifyKind1 (EUnifyKind1(..), mkEUnifyKind1) where

-- import Int

struct  Mystruct z  =
                      xx ::Int 32
                      yy ::Int 32
interface EUnifyKind1 =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32


mkEUnifyKind1 :: Module EUnifyKind1
mkEUnifyKind1 =
      module

	w :: Reg (Int 32)
	w <- mkRegU

	x :: Reg (Int 32)
	x <- mkRegU

	y :: Reg (Int 32)
	y <- mkReg 0

        z :: Mystruct
        z.xx :: Reg (Int 32)

        z.yy :: Reg (Int 32)

        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
                            let
                               (x,y) = split z
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0


