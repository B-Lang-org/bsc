function a func provisos (Bits#(a,sa), Arith#(a));
    func = unpack(0) + unpack(1);
endfunction
