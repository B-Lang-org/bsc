(* synthesize *)
(* gate_input_clocks="c1, c3" *)
module sysGateInputClocks1 #(Clock c1, Clock c2, Clock c3) ();
endmodule

