package IfMultiAction(sysMultiAction, MultiAction(..)) where

import Environment

interface MultiAction =
  f :: Bool -> Bool -> Action
  reset :: Action
  print :: Action
  finish :: Action

sysMultiAction :: Module MultiAction
sysMultiAction =
  module
    r1 :: Reg (UInt 20) <- mkReg 0
    r2 :: Reg (UInt 20) <- mkReg 0
    r3 :: Reg (UInt 20) <- mkReg 0
    r4 :: Reg (UInt 20) <- mkReg 0
    r5 :: Reg (UInt 20) <- mkReg 0

    interface
      f a b = if a then
               action {r1 :=1;
                       if b then
                          r2 := 1
                       else
                          r3 := 1;
                       r4 :=1 }
              else action { r4:=2; r5:=1; if b then r2 := 1 else r3 := 1}
      reset = action {r1:=0; r2:=0; r3:=0; r4:=0; r5:=0}
      print = $display "0x%h" (pack (r5+(16*r4)+(256*r3)+(4096*r2)+(65536*r1)))
      finish = $finish 0
