function Action f();
  action
    bit [3:0] x;
    begin
      action
      endaction
    end
  endaction
endfunction
