-----------------------------------------------------------------------
-- Project: Bluespec

-- File: ERTSOutOfMemory1.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers an "out of memory" error

-- Error Message : bsc +RTS -A4G -M4G -RTS -verilog -g mkERTSOutOfMemory1 ERTSOutOfMemory1.bs
-- bsc: out of memory (requested 1048576 bytes)
-----------------------------------------------------------------------

package ERTSOutOfMemory1 (ERTSOutOfMemory1(..), mkERTSOutOfMemory1) where

-- import Int

interface ERTSOutOfMemory1 =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32

mkERTSOutOfMemory1 :: Module ERTSOutOfMemory1
mkERTSOutOfMemory1 =
    module
        x :: Reg (Int 32)
        x <- mkRegU

        y :: Reg (Int 32)
        y <- mkReg 0

        rules
          "Swap":
            when x > y, y /= 0
              ==> action
                      x := y
                      y := x

          "Subtract":
            when x <= y, y /= 0
              ==> action
                      y := y - x

        interface
            start ix iy = action
                              x := ix
                              y := iy
                          when y == 0
            result = x when y == 0


