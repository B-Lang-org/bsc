// Define a shorthand for computing the square of a numeric type
// This is used to compute the row & column lengths given the order
// of the sudoku grid, and to compute the number of cells given the
// the row/column length.
typedef TMul#(x,x) TSquare#(numeric type x);
