//500 Rules with the descendancy attribute.

package Five_Hundred_Rules;

module mkFive_Hundred_Rules();

    Reg#(Bit#(10)) count();
    mkReg#(0) count_r(count);

    Reg#(Bit#(11)) count2();
    mkReg#(0) count2_r(count2);

    (* descending_urgency = "test_rule_500, test_rule_499, test_rule_498, test_rule_497, test_rule_496, test_rule_495, test_rule_494, test_rule_493, test_rule_492,test_rule_491, test_rule_490, test_rule_489, test_rule_488, test_rule_487, test_rule_486, test_rule_485, test_rule_484, test_rule_483, test_rule_482,test_rule_481, test_rule_480, test_rule_479, test_rule_478, test_rule_477, test_rule_476, test_rule_475, test_rule_474, test_rule_473, test_rule_472,test_rule_471, test_rule_470,  test_rule_469, test_rule_468, test_rule_467, test_rule_466, test_rule_465, test_rule_464, test_rule_463, test_rule_462,test_rule_461, test_rule_460, test_rule_459, test_rule_458, test_rule_457, test_rule_456, test_rule_455, test_rule_454, test_rule_453, test_rule_452,test_rule_451, test_rule_450,  test_rule_449, test_rule_448, test_rule_447, test_rule_446, test_rule_445, test_rule_444, test_rule_443, test_rule_442,test_rule_441, test_rule_440,test_rule_439, test_rule_438, test_rule_437, test_rule_436, test_rule_435, test_rule_434, test_rule_433, test_rule_432,test_rule_431, test_rule_430,  test_rule_429, test_rule_428, test_rule_427, test_rule_426, test_rule_425, test_rule_424, test_rule_423, test_rule_422,test_rule_421, test_rule_420,test_rule_419, test_rule_418, test_rule_417, test_rule_416, test_rule_415, test_rule_414, test_rule_413, test_rule_412,test_rule_411, test_rule_410,  test_rule_409, test_rule_408, test_rule_407, test_rule_406, test_rule_405, test_rule_404, test_rule_403, test_rule_402,test_rule_401, test_rule_400, test_rule_399, test_rule_398, test_rule_397, test_rule_396, test_rule_395, test_rule_394, test_rule_393, test_rule_392,test_rule_391, test_rule_390, test_rule_389, test_rule_388, test_rule_387, test_rule_386, test_rule_385, test_rule_384, test_rule_383, test_rule_382,test_rule_381, test_rule_380, test_rule_379, test_rule_378, test_rule_377, test_rule_376, test_rule_375, test_rule_374, test_rule_373, test_rule_372,test_rule_371, test_rule_370,  test_rule_369, test_rule_368, test_rule_367, test_rule_366, test_rule_365, test_rule_364, test_rule_363, test_rule_362,test_rule_361, test_rule_360, test_rule_359, test_rule_358, test_rule_357, test_rule_356, test_rule_355, test_rule_354, test_rule_353, test_rule_352,test_rule_351, test_rule_350,  test_rule_349, test_rule_348, test_rule_347, test_rule_346, test_rule_345, test_rule_344, test_rule_343, test_rule_342,test_rule_341, test_rule_340,test_rule_339, test_rule_338, test_rule_337, test_rule_336, test_rule_335, test_rule_334, test_rule_333, test_rule_332,test_rule_331, test_rule_330,  test_rule_329, test_rule_328, test_rule_327, test_rule_326, test_rule_325, test_rule_324, test_rule_323, test_rule_322,test_rule_321, test_rule_320,test_rule_319, test_rule_318, test_rule_317, test_rule_316, test_rule_315, test_rule_314, test_rule_313, test_rule_312,test_rule_311, test_rule_310,  test_rule_309, test_rule_308, test_rule_307, test_rule_306, test_rule_305, test_rule_304, test_rule_303, test_rule_302,test_rule_301, test_rule_300,test_rule_299, test_rule_298, test_rule_297, test_rule_296, test_rule_295, test_rule_294, test_rule_293, test_rule_292,test_rule_291, test_rule_290, test_rule_289, test_rule_288, test_rule_287, test_rule_286, test_rule_285, test_rule_284, test_rule_283, test_rule_282,test_rule_281, test_rule_280, test_rule_279, test_rule_278, test_rule_277, test_rule_276, test_rule_275, test_rule_274, test_rule_273, test_rule_272,test_rule_271, test_rule_270,  test_rule_269, test_rule_268, test_rule_267, test_rule_266, test_rule_265, test_rule_264, test_rule_263, test_rule_262,test_rule_261, test_rule_260, test_rule_259, test_rule_258, test_rule_257, test_rule_256, test_rule_255, test_rule_254, test_rule_253, test_rule_252,test_rule_251, test_rule_250,  test_rule_249, test_rule_248, test_rule_247, test_rule_246, test_rule_245, test_rule_244, test_rule_243, test_rule_242,test_rule_241, test_rule_240,test_rule_239, test_rule_238, test_rule_237, test_rule_236, test_rule_235, test_rule_234, test_rule_233, test_rule_232,test_rule_231, test_rule_230,  test_rule_229, test_rule_228, test_rule_227, test_rule_226, test_rule_225, test_rule_224, test_rule_223, test_rule_222,test_rule_221, test_rule_220,test_rule_219, test_rule_218, test_rule_217, test_rule_216, test_rule_215, test_rule_214, test_rule_213, test_rule_212,test_rule_211, test_rule_210,  test_rule_209, test_rule_208, test_rule_207, test_rule_206, test_rule_205, test_rule_204, test_rule_203, test_rule_202,test_rule_201, test_rule_200, test_rule_199, test_rule_198, test_rule_197, test_rule_196, test_rule_195, test_rule_194, test_rule_193, test_rule_192,test_rule_191, test_rule_190, test_rule_189, test_rule_188, test_rule_187, test_rule_186, test_rule_185, test_rule_184, test_rule_183, test_rule_182,test_rule_181, test_rule_180, test_rule_179, test_rule_178, test_rule_177, test_rule_176, test_rule_175, test_rule_174, test_rule_173, test_rule_172,test_rule_171, test_rule_170,  test_rule_169, test_rule_168, test_rule_167, test_rule_166, test_rule_165, test_rule_164, test_rule_163, test_rule_162,test_rule_161, test_rule_160, test_rule_159, test_rule_158, test_rule_157, test_rule_156, test_rule_155, test_rule_154, test_rule_153, test_rule_152,test_rule_151, test_rule_150,  test_rule_149, test_rule_148, test_rule_147, test_rule_146, test_rule_145, test_rule_144, test_rule_143, test_rule_142,test_rule_141, test_rule_140,test_rule_139, test_rule_138, test_rule_137, test_rule_136, test_rule_135, test_rule_134, test_rule_133, test_rule_132,test_rule_131, test_rule_130,  test_rule_129, test_rule_128, test_rule_127, test_rule_126, test_rule_125, test_rule_124, test_rule_123, test_rule_122,test_rule_121, test_rule_120,test_rule_119, test_rule_118, test_rule_117, test_rule_116, test_rule_115, test_rule_114, test_rule_113, test_rule_112,test_rule_111, test_rule_110,  test_rule_109, test_rule_108, test_rule_107, test_rule_106, test_rule_105, test_rule_104, test_rule_103, test_rule_102,test_rule_101, test_rule_100, test_rule_99, test_rule_98, test_rule_97, test_rule_96, test_rule_95, test_rule_94, test_rule_93, test_rule_92,test_rule_91, test_rule_90, test_rule_89, test_rule_88, test_rule_87, test_rule_86, test_rule_85, test_rule_84, test_rule_83, test_rule_82,test_rule_81, test_rule_80, test_rule_79, test_rule_78, test_rule_77, test_rule_76, test_rule_75, test_rule_74, test_rule_73, test_rule_72,test_rule_71, test_rule_70,  test_rule_69, test_rule_68, test_rule_67, test_rule_66, test_rule_65, test_rule_64, test_rule_63, test_rule_62,test_rule_61, test_rule_60, test_rule_59, test_rule_58, test_rule_57, test_rule_56, test_rule_55, test_rule_54, test_rule_53, test_rule_52,test_rule_51, test_rule_50,  test_rule_49, test_rule_48, test_rule_47, test_rule_46, test_rule_45, test_rule_44, test_rule_43, test_rule_42,test_rule_41, test_rule_40,test_rule_39, test_rule_38, test_rule_37, test_rule_36, test_rule_35, test_rule_34, test_rule_33, test_rule_32,test_rule_31, test_rule_30,  test_rule_29, test_rule_28, test_rule_27, test_rule_26, test_rule_25, test_rule_24, test_rule_23, test_rule_22,test_rule_21, test_rule_20,test_rule_19, test_rule_18, test_rule_17, test_rule_16, test_rule_15, test_rule_14, test_rule_13, test_rule_12,test_rule_11, test_rule_10,  test_rule_09, test_rule_08, test_rule_07, test_rule_06, test_rule_05, test_rule_04, test_rule_03, test_rule_02,test_rule_01" *)



    rule test_rule_01 (count >= 1);
        count <= count + 1;
        $display ("Executing Rule1");
    endrule

    rule test_rule_02 (count >= 2);
        count <= count + 2;
        $display ("Executing Rule2");
    endrule

    rule test_rule_03 (count >= 3);
        count <= count + 3;
        $display ("Executing Rule3");
    endrule

    rule test_rule_04 (count >= 4);
        count <= count + 4;
        $display ("Executing Rule4");
    endrule

    rule test_rule_05 (count >= 5);
        count <= count + 5;
        $display ("Executing Rule5");
    endrule

    rule test_rule_06 (count >= 6);
        count <= count + 6;
        $display ("Executing Rule6");
    endrule

    rule test_rule_07 (count >= 7);
        count <= count + 7;
        $display ("Executing Rule7");
    endrule

    rule test_rule_08 (count >= 8);
        count <= count + 8;
        $display ("Executing Rule8");
    endrule

    rule test_rule_09 (count >= 9);
        count <= count + 9;
        $display ("Executing Rule9");
    endrule

    rule test_rule_10 (count >= 10);
        count <= count + 10;
        $display ("Executing Rule10");
    endrule

    rule test_rule_11 (count >= 11);
        count <= count + 11;
        $display ("Executing Rule11");
    endrule

    rule test_rule_12 (count >= 12);
        count <= count + 12;
        $display ("Executing Rule12");
    endrule

    rule test_rule_13 (count >= 13);
        count <= count + 13;
        $display ("Executing Rule13");
    endrule

    rule test_rule_14 (count >= 14);
        count <= count + 14;
        $display ("Executing Rule14");
    endrule

    rule test_rule_15 (count >= 15);
        count <= count + 15;
        $display ("Executing Rule15");
    endrule

    rule test_rule_16 (count >= 16);
        count <= count + 16;
        $display ("Executing Rule16");
    endrule

    rule test_rule_17 (count >= 17);
        count <= count + 17;
        $display ("Executing Rule17");
    endrule

    rule test_rule_18 (count >= 18);
        count <= count + 18;
        $display ("Executing Rule18");
    endrule

    rule test_rule_19 (count >= 19);
        count <= count + 19;
        $display ("Executing Rule19");
    endrule

    rule test_rule_20 (count >= 20);
        count <= count + 20;
        $display ("Executing Rule20");
    endrule

    rule test_rule_21 (count >= 21);
        count <= count + 21;
        $display ("Executing Rule21");
    endrule

    rule test_rule_22 (count >= 22);
        count <= count + 22;
        $display ("Executing Rule22");
    endrule

    rule test_rule_23 (count >= 23);
        count <= count + 23;
        $display ("Executing Rule23");
    endrule

    rule test_rule_24 (count >= 24);
        count <= count + 24;
        $display ("Executing Rule24");
    endrule

    rule test_rule_25 (count >= 25);
        count <= count + 25;
        $display ("Executing Rule25");
    endrule

    rule test_rule_26 (count >= 26);
        count <= count + 26;
        $display ("Executing Rule26");
    endrule

    rule test_rule_27 (count >= 27);
        count <= count + 27;
        $display ("Executing Rule27");
    endrule

    rule test_rule_28 (count >= 28);
        count <= count + 28;
        $display ("Executing Rule28");
    endrule

    rule test_rule_29 (count >= 29);
        count <= count + 29;
        $display ("Executing Rule29");
    endrule

    rule test_rule_30 (count >= 30);
        count <= count + 30;
        $display ("Executing Rule30");
    endrule

    rule test_rule_31 (count >= 31);
        count <= count + 31;
        $display ("Executing Rule31");
    endrule

    rule test_rule_32 (count >= 32);
        count <= count + 32;
        $display ("Executing Rule32");
    endrule

    rule test_rule_33 (count >= 33);
        count <= count + 33;
        $display ("Executing Rule33");
    endrule

    rule test_rule_34 (count >= 34);
        count <= count + 34;
        $display ("Executing Rule34");
    endrule

    rule test_rule_35 (count >= 35);
        count <= count + 35;
        $display ("Executing Rule35");
    endrule

    rule test_rule_36 (count >= 36);
        count <= count + 36;
        $display ("Executing Rule36");
    endrule

    rule test_rule_37 (count >= 37);
        count <= count + 37;
        $display ("Executing Rule37");
    endrule

    rule test_rule_38 (count >= 38);
        count <= count + 38;
        $display ("Executing Rule38");
    endrule

    rule test_rule_39 (count >= 39);
        count <= count + 39;
        $display ("Executing Rule39");
    endrule


    rule test_rule_40 (count >= 40);
        count <= count + 40;
        $display ("Executing Rule40");
    endrule

    rule test_rule_41 (count >= 41);
        count <= count + 41;
        $display ("Executing Rule41");
    endrule

    rule test_rule_42 (count >= 42);
        count <= count + 42;
        $display ("Executing Rule42");
    endrule

    rule test_rule_43 (count >= 43);
        count <= count + 43;
        $display ("Executing Rule43");
    endrule

    rule test_rule_44 (count >= 44);
        count <= count + 44;
        $display ("Executing Rule44");
    endrule

    rule test_rule_45 (count >= 45);
        count <= count + 45;
        $display ("Executing Rule45");
    endrule

    rule test_rule_46 (count >= 46);
        count <= count + 46;
        $display ("Executing Rule46");
    endrule

    rule test_rule_47 (count >= 47);
        count <= count + 47;
        $display ("Executing Rule47");
    endrule

    rule test_rule_48 (count >= 48);
        count <= count + 48;
        $display ("Executing Rule48");
    endrule

    rule test_rule_49 (count >= 49);
        count <= count + 49;
        $display ("Executing Rule49");
    endrule


    rule test_rule_50 (count >= 50);
        count <= count + 50;
        $display ("Executing Rule50");
    endrule

    rule test_rule_51 (count >= 51);
        count <= count + 51;
        $display ("Executing Rule51");
    endrule

    rule test_rule_52 (count >= 52);
        count <= count + 52;
        $display ("Executing Rule52");
    endrule

    rule test_rule_53 (count >= 53);
        count <= count + 53;
        $display ("Executing Rule53");
    endrule

    rule test_rule_54 (count >= 54);
        count <= count + 54;
        $display ("Executing Rule54");
    endrule

    rule test_rule_55 (count >= 55);
        count <= count + 55;
        $display ("Executing Rule55");
    endrule

    rule test_rule_56 (count >= 56);
        count <= count + 56;
        $display ("Executing Rule56");
    endrule

    rule test_rule_57 (count >= 57);
        count <= count + 57;
        $display ("Executing Rule57");
    endrule

    rule test_rule_58 (count >= 58);
        count <= count + 58;
        $display ("Executing Rule58");
    endrule

    rule test_rule_59 (count >= 59);
        count <= count + 59;
        $display ("Executing Rule59");
    endrule


    rule test_rule_60 (count >= 60);
        count <= count + 60;
        $display ("Executing Rule60");
    endrule

    rule test_rule_61 (count >= 61);
        count <= count + 61;
        $display ("Executing Rule61");
    endrule

    rule test_rule_62 (count >= 62);
        count <= count + 62;
        $display ("Executing Rule62");
    endrule

    rule test_rule_63 (count >= 63);
        count <= count + 63;
        $display ("Executing Rule63");
    endrule

    rule test_rule_64 (count >= 64);
        count <= count + 64;
        $display ("Executing Rule64");
    endrule

    rule test_rule_65 (count >= 65);
        count <= count + 65;
        $display ("Executing Rule65");
    endrule

    rule test_rule_66 (count >= 66);
        count <= count + 66;
        $display ("Executing Rule66");
    endrule

    rule test_rule_67 (count >= 67);
        count <= count + 67;
        $display ("Executing Rule67");
    endrule

    rule test_rule_68 (count >= 68);
        count <= count + 68;
        $display ("Executing Rule68");
    endrule

    rule test_rule_69 (count >= 69);
        count <= count + 69;
        $display ("Executing Rule69");
    endrule


    rule test_rule_70 (count >= 70);
        count <= count + 70;
        $display ("Executing Rule70");
    endrule

    rule test_rule_71 (count >= 71);
        count <= count + 71;
        $display ("Executing Rule71");
    endrule

    rule test_rule_72 (count >= 72);
        count <= count + 72;
        $display ("Executing Rule72");
    endrule

    rule test_rule_73 (count >= 73);
        count <= count + 73;
        $display ("Executing Rule73");
    endrule

    rule test_rule_74 (count >= 74);
        count <= count + 74;
        $display ("Executing Rule74");
    endrule

    rule test_rule_75 (count >= 75);
        count <= count + 75;
        $display ("Executing Rule75");
    endrule

    rule test_rule_76 (count >= 76);
        count <= count + 76;
        $display ("Executing Rule76");
    endrule

    rule test_rule_77 (count >= 77);
        count <= count + 77;
        $display ("Executing Rule77");
    endrule

    rule test_rule_78 (count >= 78);
        count <= count + 78;
        $display ("Executing Rule78");
    endrule

    rule test_rule_79 (count >= 79);
        count <= count + 79;
        $display ("Executing Rule79");
    endrule


    rule test_rule_80 (count >= 80);
        count <= count + 80;
        $display ("Executing Rule80");
    endrule

    rule test_rule_81 (count >= 81);
        count <= count + 81;
        $display ("Executing Rule81");
    endrule

    rule test_rule_82 (count >= 82);
        count <= count + 82;
        $display ("Executing Rule82");
    endrule

    rule test_rule_83 (count >= 83);
        count <= count + 83;
        $display ("Executing Rule83");
    endrule

    rule test_rule_84 (count >= 84);
        count <= count + 84;
        $display ("Executing Rule84");
    endrule

    rule test_rule_85 (count >= 85);
        count <= count + 85;
        $display ("Executing Rule85");
    endrule

    rule test_rule_86 (count >= 86);
        count <= count + 86;
        $display ("Executing Rule86");
    endrule

    rule test_rule_87 (count >= 87);
        count <= count + 87;
        $display ("Executing Rule87");
    endrule

    rule test_rule_88 (count >= 88);
        count <= count + 88;
        $display ("Executing Rule88");
    endrule

    rule test_rule_89 (count >= 89);
        count <= count + 89;
        $display ("Executing Rule89");
    endrule


    rule test_rule_90 (count >= 90);
        count <= count + 90;
        $display ("Executing Rule90");
    endrule

    rule test_rule_91 (count >= 91);
        count <= count + 91;
        $display ("Executing Rule91");
    endrule

    rule test_rule_92 (count >= 92);
        count <= count + 92;
        $display ("Executing Rule92");
    endrule

    rule test_rule_93 (count >= 93);
        count <= count + 93;
        $display ("Executing Rule93");
    endrule

    rule test_rule_94 (count >= 94);
        count <= count + 94;
        $display ("Executing Rule94");
    endrule

    rule test_rule_95 (count >= 95);
        count <= count + 95;
        $display ("Executing Rule95");
    endrule

    rule test_rule_96 (count >= 96);
        count <= count + 96;
        $display ("Executing Rule96");
    endrule

    rule test_rule_97 (count >= 97);
        count <= count + 97;
        $display ("Executing Rule97");
    endrule

    rule test_rule_98 (count >= 98);
        count <= count + 98;
        $display ("Executing Rule98");
    endrule

    rule test_rule_99 (count >= 99);
        count <= count + 99;
        $display ("Executing Rule99");
    endrule

    rule test_rule_100 (count >= 100);
        count <= count + 100;
        $display ("Executing Rule100");
    endrule

    rule test_rule_101 (count >= 101);
        count <= count + 101;
        $display ("Executing Rule101");
    endrule

    rule test_rule_102 (count >= 102);
        count <= count + 102;
        $display ("Executing Rule102");
    endrule

    rule test_rule_103 (count >= 103);
        count <= count + 103;
        $display ("Executing Rule103");
    endrule

    rule test_rule_104 (count >= 104);
        count <= count + 104;
        $display ("Executing Rule104");
    endrule

    rule test_rule_105 (count >= 105);
        count <= count + 105;
        $display ("Executing Rule105");
    endrule

    rule test_rule_106 (count >= 106);
        count <= count + 106;
        $display ("Executing Rule106");
    endrule

    rule test_rule_107 (count >= 107);
        count <= count + 107;
        $display ("Executing Rule107");
    endrule

    rule test_rule_108 (count >= 108);
        count <= count + 108;
        $display ("Executing Rule108");
    endrule

    rule test_rule_109 (count >= 109);
        count <= count + 109;
        $display ("Executing Rule109");
    endrule

    rule test_rule_110 (count >= 110);
        count <= count + 110;
        $display ("Executing Rule110");
    endrule

    rule test_rule_111 (count >= 111);
        count <= count + 111;
        $display ("Executing Rule111");
    endrule

    rule test_rule_112 (count >= 112);
        count <= count + 112;
        $display ("Executing Rule112");
    endrule

    rule test_rule_113 (count >= 113);
        count <= count + 113;
        $display ("Executing Rule113");
    endrule

    rule test_rule_114 (count >= 114);
        count <= count + 114;
        $display ("Executing Rule114");
    endrule

    rule test_rule_115 (count >= 115);
        count <= count + 115;
        $display ("Executing Rule115");
    endrule

    rule test_rule_116 (count >= 116);
        count <= count + 116;
        $display ("Executing Rule116");
    endrule

    rule test_rule_117 (count >= 117);
        count <= count + 117;
        $display ("Executing Rule117");
    endrule

    rule test_rule_118 (count >= 118);
        count <= count + 118;
        $display ("Executing Rule118");
    endrule

    rule test_rule_119 (count >= 119);
        count <= count + 119;
        $display ("Executing Rule119");
    endrule

    rule test_rule_120 (count >= 120);
        count <= count + 120;
        $display ("Executing Rule120");
    endrule

    rule test_rule_121 (count >= 121);
        count <= count + 121;
        $display ("Executing Rule121");
    endrule

    rule test_rule_122 (count >= 122);
        count <= count + 122;
        $display ("Executing Rule122");
    endrule

    rule test_rule_123 (count >= 123);
        count <= count + 123;
        $display ("Executing Rule123");
    endrule

    rule test_rule_124 (count >= 124);
        count <= count + 124;
        $display ("Executing Rule124");
    endrule

    rule test_rule_125 (count >= 125);
        count <= count + 125;
        $display ("Executing Rule125");
    endrule

    rule test_rule_126 (count >= 126);
        count <= count + 126;
        $display ("Executing Rule126");
    endrule

    rule test_rule_127 (count >= 127);
        count <= count + 127;
        $display ("Executing Rule127");
    endrule

    rule test_rule_128 (count >= 128);
        count <= count + 128;
        $display ("Executing Rule128");
    endrule

    rule test_rule_129 (count >= 129);
        count <= count + 129;
        $display ("Executing Rule129");
    endrule

    rule test_rule_130 (count >= 130);
        count <= count + 130;
        $display ("Executing Rule130");
    endrule

    rule test_rule_131 (count >= 131);
        count <= count + 131;
        $display ("Executing Rule131");
    endrule

    rule test_rule_132 (count >= 132);
        count <= count + 132;
        $display ("Executing Rule132");
    endrule

    rule test_rule_133 (count >= 133);
        count <= count + 133;
        $display ("Executing Rule133");
    endrule

    rule test_rule_134 (count >= 134);
        count <= count + 134;
        $display ("Executing Rule134");
    endrule

    rule test_rule_135 (count >= 135);
        count <= count + 135;
        $display ("Executing Rule135");
    endrule

    rule test_rule_136 (count >= 136);
        count <= count + 136;
        $display ("Executing Rule136");
    endrule

    rule test_rule_137 (count >= 137);
        count <= count + 137;
        $display ("Executing Rule137");
    endrule

    rule test_rule_138 (count >= 138);
        count <= count + 138;
        $display ("Executing Rule138");
    endrule

    rule test_rule_139 (count >= 139);
        count <= count + 139;
        $display ("Executing Rule139");
    endrule


    rule test_rule_140 (count >= 140);
        count <= count + 140;
        $display ("Executing Rule140");
    endrule

    rule test_rule_141 (count >= 141);
        count <= count + 141;
        $display ("Executing Rule141");
    endrule

    rule test_rule_142 (count >= 142);
        count <= count + 142;
        $display ("Executing Rule142");
    endrule

    rule test_rule_143 (count >= 143);
        count <= count + 143;
        $display ("Executing Rule143");
    endrule

    rule test_rule_144 (count >= 144);
        count <= count + 144;
        $display ("Executing Rule144");
    endrule

    rule test_rule_145 (count >= 145);
        count <= count + 145;
        $display ("Executing Rule145");
    endrule

    rule test_rule_146 (count >= 146);
        count <= count + 146;
        $display ("Executing Rule146");
    endrule

    rule test_rule_147 (count >= 147);
        count <= count + 147;
        $display ("Executing Rule147");
    endrule

    rule test_rule_148 (count >= 148);
        count <= count + 148;
        $display ("Executing Rule148");
    endrule

    rule test_rule_149 (count >= 149);
        count <= count + 149;
        $display ("Executing Rule149");
    endrule


    rule test_rule_150 (count >= 150);
        count <= count + 150;
        $display ("Executing Rule150");
    endrule

    rule test_rule_151 (count >= 151);
        count <= count + 151;
        $display ("Executing Rule151");
    endrule

    rule test_rule_152 (count >= 152);
        count <= count + 152;
        $display ("Executing Rule152");
    endrule

    rule test_rule_153 (count >= 153);
        count <= count + 153;
        $display ("Executing Rule153");
    endrule

    rule test_rule_154 (count >= 154);
        count <= count + 154;
        $display ("Executing Rule154");
    endrule

    rule test_rule_155 (count >= 155);
        count <= count + 155;
        $display ("Executing Rule155");
    endrule

    rule test_rule_156 (count >= 156);
        count <= count + 156;
        $display ("Executing Rule156");
    endrule

    rule test_rule_157 (count >= 157);
        count <= count + 157;
        $display ("Executing Rule157");
    endrule

    rule test_rule_158 (count >= 158);
        count <= count + 158;
        $display ("Executing Rule158");
    endrule

    rule test_rule_159 (count >= 159);
        count <= count + 159;
        $display ("Executing Rule159");
    endrule


    rule test_rule_160 (count >= 160);
        count <= count + 160;
        $display ("Executing Rule160");
    endrule

    rule test_rule_161 (count >= 161);
        count <= count + 161;
        $display ("Executing Rule161");
    endrule

    rule test_rule_162 (count >= 162);
        count <= count + 162;
        $display ("Executing Rule162");
    endrule

    rule test_rule_163 (count >= 163);
        count <= count + 163;
        $display ("Executing Rule163");
    endrule

    rule test_rule_164 (count >= 164);
        count <= count + 164;
        $display ("Executing Rule164");
    endrule

    rule test_rule_165 (count >= 165);
        count <= count + 165;
        $display ("Executing Rule165");
    endrule

    rule test_rule_166 (count >= 166);
        count <= count + 166;
        $display ("Executing Rule166");
    endrule

    rule test_rule_167 (count >= 167);
        count <= count + 167;
        $display ("Executing Rule167");
    endrule

    rule test_rule_168 (count >= 168);
        count <= count + 168;
        $display ("Executing Rule168");
    endrule

    rule test_rule_169 (count >= 169);
        count <= count + 169;
        $display ("Executing Rule169");
    endrule


    rule test_rule_170 (count >= 170);
        count <= count + 170;
        $display ("Executing Rule170");
    endrule

    rule test_rule_171 (count >= 171);
        count <= count + 171;
        $display ("Executing Rule171");
    endrule

    rule test_rule_172 (count >= 172);
        count <= count + 172;
        $display ("Executing Rule172");
    endrule

    rule test_rule_173 (count >= 173);
        count <= count + 173;
        $display ("Executing Rule173");
    endrule

    rule test_rule_174 (count >= 174);
        count <= count + 174;
        $display ("Executing Rule174");
    endrule

    rule test_rule_175 (count >= 175);
        count <= count + 175;
        $display ("Executing Rule175");
    endrule

    rule test_rule_176 (count >= 176);
        count <= count + 176;
        $display ("Executing Rule176");
    endrule

    rule test_rule_177 (count >= 177);
        count <= count + 177;
        $display ("Executing Rule177");
    endrule

    rule test_rule_178 (count >= 178);
        count <= count + 178;
        $display ("Executing Rule178");
    endrule

    rule test_rule_179 (count >= 179);
        count <= count + 179;
        $display ("Executing Rule179");
    endrule


    rule test_rule_180 (count >= 180);
        count <= count + 180;
        $display ("Executing Rule180");
    endrule

    rule test_rule_181 (count >= 181);
        count <= count + 181;
        $display ("Executing Rule181");
    endrule

    rule test_rule_182 (count >= 182);
        count <= count + 182;
        $display ("Executing Rule182");
    endrule

    rule test_rule_183 (count >= 183);
        count <= count + 183;
        $display ("Executing Rule183");
    endrule

    rule test_rule_184 (count >= 184);
        count <= count + 184;
        $display ("Executing Rule184");
    endrule

    rule test_rule_185 (count >= 185);
        count <= count + 185;
        $display ("Executing Rule185");
    endrule

    rule test_rule_186 (count >= 186);
        count <= count + 186;
        $display ("Executing Rule186");
    endrule

    rule test_rule_187 (count >= 187);
        count <= count + 187;
        $display ("Executing Rule187");
    endrule

    rule test_rule_188 (count >= 188);
        count <= count + 188;
        $display ("Executing Rule188");
    endrule

    rule test_rule_189 (count >= 189);
        count <= count + 189;
        $display ("Executing Rule189");
    endrule


    rule test_rule_190 (count >= 190);
        count <= count + 190;
        $display ("Executing Rule190");
    endrule

    rule test_rule_191 (count >= 191);
        count <= count + 191;
        $display ("Executing Rule191");
    endrule

    rule test_rule_192 (count >= 192);
        count <= count + 192;
        $display ("Executing Rule192");
    endrule

    rule test_rule_193 (count >= 193);
        count <= count + 193;
        $display ("Executing Rule193");
    endrule

    rule test_rule_194 (count >= 194);
        count <= count + 194;
        $display ("Executing Rule194");
    endrule

    rule test_rule_195 (count >= 195);
        count <= count + 195;
        $display ("Executing Rule195");
    endrule

    rule test_rule_196 (count >= 196);
        count <= count + 196;
        $display ("Executing Rule196");
    endrule

    rule test_rule_197 (count >= 197);
        count <= count + 197;
        $display ("Executing Rule197");
    endrule

    rule test_rule_198 (count >= 198);
        count <= count + 198;
        $display ("Executing Rule198");
    endrule

    rule test_rule_199 (count >= 199);
        count <= count + 199;
        $display ("Executing Rule199");
    endrule




    rule test_rule_200 (count >= 200);
        count <= count + 200;
        $display ("Executing Rule200");
    endrule

    rule test_rule_201 (count >= 201);
        count <= count + 201;
        $display ("Executing Rule201");
    endrule

    rule test_rule_202 (count >= 202);
        count <= count + 202;
        $display ("Executing Rule202");
    endrule

    rule test_rule_203 (count >= 203);
        count <= count + 203;
        $display ("Executing Rule203");
    endrule

    rule test_rule_204 (count >= 204);
        count <= count + 204;
        $display ("Executing Rule204");
    endrule

    rule test_rule_205 (count >= 205);
        count <= count + 205;
        $display ("Executing Rule205");
    endrule

    rule test_rule_206 (count >= 206);
        count <= count + 206;
        $display ("Executing Rule206");
    endrule

    rule test_rule_207 (count >= 207);
        count <= count + 207;
        $display ("Executing Rule207");
    endrule

    rule test_rule_208 (count >= 208);
        count <= count + 208;
        $display ("Executing Rule208");
    endrule

    rule test_rule_209 (count >= 209);
        count <= count + 209;
        $display ("Executing Rule209");
    endrule

    rule test_rule_210 (count >= 210);
        count <= count + 210;
        $display ("Executing Rule210");
    endrule

    rule test_rule_211 (count >= 211);
        count <= count + 211;
        $display ("Executing Rule211");
    endrule

    rule test_rule_212 (count >= 212);
        count <= count + 212;
        $display ("Executing Rule212");
    endrule

    rule test_rule_213 (count >= 213);
        count <= count + 213;
        $display ("Executing Rule213");
    endrule

    rule test_rule_214 (count >= 214);
        count <= count + 214;
        $display ("Executing Rule214");
    endrule

    rule test_rule_215 (count >= 215);
        count <= count + 215;
        $display ("Executing Rule215");
    endrule

    rule test_rule_216 (count >= 216);
        count <= count + 216;
        $display ("Executing Rule216");
    endrule

    rule test_rule_217 (count >= 217);
        count <= count + 217;
        $display ("Executing Rule217");
    endrule

    rule test_rule_218 (count >= 218);
        count <= count + 218;
        $display ("Executing Rule218");
    endrule

    rule test_rule_219 (count >= 219);
        count <= count + 219;
        $display ("Executing Rule219");
    endrule

    rule test_rule_220 (count >= 220);
        count <= count + 220;
        $display ("Executing Rule220");
    endrule

    rule test_rule_221 (count >= 221);
        count <= count + 221;
        $display ("Executing Rule221");
    endrule

    rule test_rule_222 (count >= 222);
        count <= count + 222;
        $display ("Executing Rule222");
    endrule

    rule test_rule_223 (count >= 223);
        count <= count + 223;
        $display ("Executing Rule223");
    endrule

    rule test_rule_224 (count >= 224);
        count <= count + 224;
        $display ("Executing Rule224");
    endrule

    rule test_rule_225 (count >= 225);
        count <= count + 225;
        $display ("Executing Rule225");
    endrule

    rule test_rule_226 (count >= 226);
        count <= count + 226;
        $display ("Executing Rule226");
    endrule

    rule test_rule_227 (count >= 227);
        count <= count + 227;
        $display ("Executing Rule227");
    endrule

    rule test_rule_228 (count >= 228);
        count <= count + 228;
        $display ("Executing Rule228");
    endrule

    rule test_rule_229 (count >= 229);
        count <= count + 229;
        $display ("Executing Rule229");
    endrule

    rule test_rule_230 (count >= 230);
        count <= count + 230;
        $display ("Executing Rule230");
    endrule

    rule test_rule_231 (count >= 231);
        count <= count + 231;
        $display ("Executing Rule231");
    endrule

    rule test_rule_232 (count >= 232);
        count <= count + 232;
        $display ("Executing Rule232");
    endrule

    rule test_rule_233 (count >= 233);
        count <= count + 233;
        $display ("Executing Rule233");
    endrule

    rule test_rule_234 (count >= 234);
        count <= count + 234;
        $display ("Executing Rule234");
    endrule

    rule test_rule_235 (count >= 235);
        count <= count + 235;
        $display ("Executing Rule235");
    endrule

    rule test_rule_236 (count >= 236);
        count <= count + 236;
        $display ("Executing Rule236");
    endrule

    rule test_rule_237 (count >= 237);
        count <= count + 237;
        $display ("Executing Rule237");
    endrule

    rule test_rule_238 (count >= 238);
        count <= count + 238;
        $display ("Executing Rule238");
    endrule

    rule test_rule_239 (count >= 239);
        count <= count + 239;
        $display ("Executing Rule239");
    endrule


    rule test_rule_240 (count >= 240);
        count <= count + 240;
        $display ("Executing Rule240");
    endrule

    rule test_rule_241 (count >= 241);
        count <= count + 241;
        $display ("Executing Rule241");
    endrule

    rule test_rule_242 (count >= 242);
        count <= count + 242;
        $display ("Executing Rule242");
    endrule

    rule test_rule_243 (count >= 243);
        count <= count + 243;
        $display ("Executing Rule243");
    endrule

    rule test_rule_244 (count >= 244);
        count <= count + 244;
        $display ("Executing Rule244");
    endrule

    rule test_rule_245 (count >= 245);
        count <= count + 245;
        $display ("Executing Rule245");
    endrule

    rule test_rule_246 (count >= 246);
        count <= count + 246;
        $display ("Executing Rule246");
    endrule

    rule test_rule_247 (count >= 247);
        count <= count + 247;
        $display ("Executing Rule247");
    endrule

    rule test_rule_248 (count >= 248);
        count <= count + 248;
        $display ("Executing Rule248");
    endrule

    rule test_rule_249 (count >= 249);
        count <= count + 249;
        $display ("Executing Rule249");
    endrule


    rule test_rule_250 (count >= 250);
        count <= count + 250;
        $display ("Executing Rule250");
    endrule

    rule test_rule_251 (count >= 251);
        count <= count + 251;
        $display ("Executing Rule251");
    endrule

    rule test_rule_252 (count >= 252);
        count <= count + 252;
        $display ("Executing Rule252");
    endrule

    rule test_rule_253 (count >= 253);
        count <= count + 253;
        $display ("Executing Rule253");
    endrule

    rule test_rule_254 (count >= 254);
        count <= count + 254;
        $display ("Executing Rule254");
    endrule

    rule test_rule_255 (count >= 255);
        count <= count + 255;
        $display ("Executing Rule255");
    endrule

    rule test_rule_256 (count >= 256);
        count <= count + 256;
        $display ("Executing Rule256");
    endrule

    rule test_rule_257 (count >= 257);
        count <= count + 257;
        $display ("Executing Rule257");
    endrule

    rule test_rule_258 (count >= 258);
        count <= count + 258;
        $display ("Executing Rule258");
    endrule

    rule test_rule_259 (count >= 259);
        count <= count + 259;
        $display ("Executing Rule259");
    endrule


    rule test_rule_260 (count >= 260);
        count <= count + 260;
        $display ("Executing Rule260");
    endrule

    rule test_rule_261 (count >= 261);
        count <= count + 261;
        $display ("Executing Rule261");
    endrule

    rule test_rule_262 (count >= 262);
        count <= count + 262;
        $display ("Executing Rule262");
    endrule

    rule test_rule_263 (count >= 263);
        count <= count + 263;
        $display ("Executing Rule263");
    endrule

    rule test_rule_264 (count >= 264);
        count <= count + 264;
        $display ("Executing Rule264");
    endrule

    rule test_rule_265 (count >= 265);
        count <= count + 265;
        $display ("Executing Rule265");
    endrule

    rule test_rule_266 (count >= 266);
        count <= count + 266;
        $display ("Executing Rule266");
    endrule

    rule test_rule_267 (count >= 267);
        count <= count + 267;
        $display ("Executing Rule267");
    endrule

    rule test_rule_268 (count >= 268);
        count <= count + 268;
        $display ("Executing Rule268");
    endrule

    rule test_rule_269 (count >= 269);
        count <= count + 269;
        $display ("Executing Rule269");
    endrule


    rule test_rule_270 (count >= 270);
        count <= count + 270;
        $display ("Executing Rule270");
    endrule

    rule test_rule_271 (count >= 271);
        count <= count + 271;
        $display ("Executing Rule271");
    endrule

    rule test_rule_272 (count >= 272);
        count <= count + 272;
        $display ("Executing Rule272");
    endrule

    rule test_rule_273 (count >= 273);
        count <= count + 273;
        $display ("Executing Rule273");
    endrule

    rule test_rule_274 (count >= 274);
        count <= count + 274;
        $display ("Executing Rule274");
    endrule

    rule test_rule_275 (count >= 275);
        count <= count + 275;
        $display ("Executing Rule275");
    endrule

    rule test_rule_276 (count >= 276);
        count <= count + 276;
        $display ("Executing Rule276");
    endrule

    rule test_rule_277 (count >= 277);
        count <= count + 277;
        $display ("Executing Rule277");
    endrule

    rule test_rule_278 (count >= 278);
        count <= count + 278;
        $display ("Executing Rule278");
    endrule

    rule test_rule_279 (count >= 279);
        count <= count + 279;
        $display ("Executing Rule279");
    endrule


    rule test_rule_280 (count >= 280);
        count <= count + 280;
        $display ("Executing Rule280");
    endrule

    rule test_rule_281 (count >= 281);
        count <= count + 281;
        $display ("Executing Rule281");
    endrule

    rule test_rule_282 (count >= 282);
        count <= count + 282;
        $display ("Executing Rule282");
    endrule

    rule test_rule_283 (count >= 283);
        count <= count + 283;
        $display ("Executing Rule283");
    endrule

    rule test_rule_284 (count >= 284);
        count <= count + 284;
        $display ("Executing Rule284");
    endrule

    rule test_rule_285 (count >= 285);
        count <= count + 285;
        $display ("Executing Rule285");
    endrule

    rule test_rule_286 (count >= 286);
        count <= count + 286;
        $display ("Executing Rule286");
    endrule

    rule test_rule_287 (count >= 287);
        count <= count + 287;
        $display ("Executing Rule287");
    endrule

    rule test_rule_288 (count >= 288);
        count <= count + 288;
        $display ("Executing Rule288");
    endrule

    rule test_rule_289 (count >= 289);
        count <= count + 289;
        $display ("Executing Rule289");
    endrule


    rule test_rule_290 (count >= 290);
        count <= count + 290;
        $display ("Executing Rule290");
    endrule

    rule test_rule_291 (count >= 291);
        count <= count + 291;
        $display ("Executing Rule291");
    endrule

    rule test_rule_292 (count >= 292);
        count <= count + 292;
        $display ("Executing Rule292");
    endrule

    rule test_rule_293 (count >= 293);
        count <= count + 293;
        $display ("Executing Rule293");
    endrule

    rule test_rule_294 (count >= 294);
        count <= count + 294;
        $display ("Executing Rule294");
    endrule

    rule test_rule_295 (count >= 295);
        count <= count + 295;
        $display ("Executing Rule295");
    endrule

    rule test_rule_296 (count >= 296);
        count <= count + 296;
        $display ("Executing Rule296");
    endrule

    rule test_rule_297 (count >= 297);
        count <= count + 297;
        $display ("Executing Rule297");
    endrule

    rule test_rule_298 (count >= 298);
        count <= count + 298;
        $display ("Executing Rule298");
    endrule

    rule test_rule_299 (count >= 299);
        count <= count + 299;
        $display ("Executing Rule299");
    endrule



    rule test_rule_300 (count >= 300);
        count <= count + 300;
        $display ("Executing Rule300");
    endrule

    rule test_rule_301 (count >= 301);
        count <= count + 301;
        $display ("Executing Rule301");
    endrule

    rule test_rule_302 (count >= 302);
        count <= count + 302;
        $display ("Executing Rule302");
    endrule

    rule test_rule_303 (count >= 303);
        count <= count + 303;
        $display ("Executing Rule303");
    endrule

    rule test_rule_304 (count >= 304);
        count <= count + 304;
        $display ("Executing Rule304");
    endrule

    rule test_rule_305 (count >= 305);
        count <= count + 305;
        $display ("Executing Rule305");
    endrule

    rule test_rule_306 (count >= 306);
        count <= count + 306;
        $display ("Executing Rule306");
    endrule

    rule test_rule_307 (count >= 307);
        count <= count + 307;
        $display ("Executing Rule307");
    endrule

    rule test_rule_308 (count >= 308);
        count <= count + 308;
        $display ("Executing Rule308");
    endrule

    rule test_rule_309 (count >= 309);
        count <= count + 309;
        $display ("Executing Rule309");
    endrule

    rule test_rule_310 (count >= 310);
        count <= count + 310;
        $display ("Executing Rule310");
    endrule

    rule test_rule_311 (count >= 311);
        count <= count + 311;
        $display ("Executing Rule311");
    endrule

    rule test_rule_312 (count >= 312);
        count <= count + 312;
        $display ("Executing Rule312");
    endrule

    rule test_rule_313 (count >= 313);
        count <= count + 313;
        $display ("Executing Rule313");
    endrule

    rule test_rule_314 (count >= 314);
        count <= count + 314;
        $display ("Executing Rule314");
    endrule

    rule test_rule_315 (count >= 315);
        count <= count + 315;
        $display ("Executing Rule315");
    endrule

    rule test_rule_316 (count >= 316);
        count <= count + 316;
        $display ("Executing Rule316");
    endrule

    rule test_rule_317 (count >= 317);
        count <= count + 317;
        $display ("Executing Rule317");
    endrule

    rule test_rule_318 (count >= 318);
        count <= count + 318;
        $display ("Executing Rule318");
    endrule

    rule test_rule_319 (count >= 319);
        count <= count + 319;
        $display ("Executing Rule319");
    endrule

    rule test_rule_320 (count >= 320);
        count <= count + 320;
        $display ("Executing Rule320");
    endrule

    rule test_rule_321 (count >= 321);
        count <= count + 321;
        $display ("Executing Rule321");
    endrule

    rule test_rule_322 (count >= 322);
        count <= count + 322;
        $display ("Executing Rule322");
    endrule

    rule test_rule_323 (count >= 323);
        count <= count + 323;
        $display ("Executing Rule323");
    endrule

    rule test_rule_324 (count >= 324);
        count <= count + 324;
        $display ("Executing Rule324");
    endrule

    rule test_rule_325 (count >= 325);
        count <= count + 325;
        $display ("Executing Rule325");
    endrule

    rule test_rule_326 (count >= 326);
        count <= count + 326;
        $display ("Executing Rule326");
    endrule

    rule test_rule_327 (count >= 327);
        count <= count + 327;
        $display ("Executing Rule327");
    endrule

    rule test_rule_328 (count >= 328);
        count <= count + 328;
        $display ("Executing Rule328");
    endrule

    rule test_rule_329 (count >= 329);
        count <= count + 329;
        $display ("Executing Rule329");
    endrule

    rule test_rule_330 (count >= 330);
        count <= count + 330;
        $display ("Executing Rule330");
    endrule

    rule test_rule_331 (count >= 331);
        count <= count + 331;
        $display ("Executing Rule331");
    endrule

    rule test_rule_332 (count >= 332);
        count <= count + 332;
        $display ("Executing Rule332");
    endrule

    rule test_rule_333 (count >= 333);
        count <= count + 333;
        $display ("Executing Rule333");
    endrule

    rule test_rule_334 (count >= 334);
        count <= count + 334;
        $display ("Executing Rule334");
    endrule

    rule test_rule_335 (count >= 335);
        count <= count + 335;
        $display ("Executing Rule335");
    endrule

    rule test_rule_336 (count >= 336);
        count <= count + 336;
        $display ("Executing Rule336");
    endrule

    rule test_rule_337 (count >= 337);
        count <= count + 337;
        $display ("Executing Rule337");
    endrule

    rule test_rule_338 (count >= 338);
        count <= count + 338;
        $display ("Executing Rule338");
    endrule

    rule test_rule_339 (count >= 339);
        count <= count + 339;
        $display ("Executing Rule339");
    endrule


    rule test_rule_340 (count >= 340);
        count <= count + 340;
        $display ("Executing Rule340");
    endrule

    rule test_rule_341 (count >= 341);
        count <= count + 341;
        $display ("Executing Rule341");
    endrule

    rule test_rule_342 (count >= 342);
        count <= count + 342;
        $display ("Executing Rule342");
    endrule

    rule test_rule_343 (count >= 343);
        count <= count + 343;
        $display ("Executing Rule343");
    endrule

    rule test_rule_344 (count >= 344);
        count <= count + 344;
        $display ("Executing Rule344");
    endrule

    rule test_rule_345 (count >= 345);
        count <= count + 345;
        $display ("Executing Rule345");
    endrule

    rule test_rule_346 (count >= 346);
        count <= count + 346;
        $display ("Executing Rule346");
    endrule

    rule test_rule_347 (count >= 347);
        count <= count + 347;
        $display ("Executing Rule347");
    endrule

    rule test_rule_348 (count >= 348);
        count <= count + 348;
        $display ("Executing Rule348");
    endrule

    rule test_rule_349 (count >= 349);
        count <= count + 349;
        $display ("Executing Rule349");
    endrule


    rule test_rule_350 (count >= 350);
        count <= count + 350;
        $display ("Executing Rule350");
    endrule

    rule test_rule_351 (count >= 351);
        count <= count + 351;
        $display ("Executing Rule351");
    endrule

    rule test_rule_352 (count >= 352);
        count <= count + 352;
        $display ("Executing Rule352");
    endrule

    rule test_rule_353 (count >= 353);
        count <= count + 353;
        $display ("Executing Rule353");
    endrule

    rule test_rule_354 (count >= 354);
        count <= count + 354;
        $display ("Executing Rule354");
    endrule

    rule test_rule_355 (count >= 355);
        count <= count + 355;
        $display ("Executing Rule355");
    endrule

    rule test_rule_356 (count >= 356);
        count <= count + 356;
        $display ("Executing Rule356");
    endrule

    rule test_rule_357 (count >= 357);
        count <= count + 357;
        $display ("Executing Rule357");
    endrule

    rule test_rule_358 (count >= 358);
        count <= count + 358;
        $display ("Executing Rule358");
    endrule

    rule test_rule_359 (count >= 359);
        count <= count + 359;
        $display ("Executing Rule359");
    endrule


    rule test_rule_360 (count >= 360);
        count <= count + 360;
        $display ("Executing Rule360");
    endrule

    rule test_rule_361 (count >= 361);
        count <= count + 361;
        $display ("Executing Rule361");
    endrule

    rule test_rule_362 (count >= 362);
        count <= count + 362;
        $display ("Executing Rule362");
    endrule

    rule test_rule_363 (count >= 363);
        count <= count + 363;
        $display ("Executing Rule363");
    endrule

    rule test_rule_364 (count >= 364);
        count <= count + 364;
        $display ("Executing Rule364");
    endrule

    rule test_rule_365 (count >= 365);
        count <= count + 365;
        $display ("Executing Rule365");
    endrule

    rule test_rule_366 (count >= 366);
        count <= count + 366;
        $display ("Executing Rule366");
    endrule

    rule test_rule_367 (count >= 367);
        count <= count + 367;
        $display ("Executing Rule367");
    endrule

    rule test_rule_368 (count >= 368);
        count <= count + 368;
        $display ("Executing Rule368");
    endrule

    rule test_rule_369 (count >= 369);
        count <= count + 369;
        $display ("Executing Rule369");
    endrule


    rule test_rule_370 (count >= 370);
        count <= count + 370;
        $display ("Executing Rule370");
    endrule

    rule test_rule_371 (count >= 371);
        count <= count + 371;
        $display ("Executing Rule371");
    endrule

    rule test_rule_372 (count >= 372);
        count <= count + 372;
        $display ("Executing Rule372");
    endrule

    rule test_rule_373 (count >= 373);
        count <= count + 373;
        $display ("Executing Rule373");
    endrule

    rule test_rule_374 (count >= 374);
        count <= count + 374;
        $display ("Executing Rule374");
    endrule

    rule test_rule_375 (count >= 375);
        count <= count + 375;
        $display ("Executing Rule375");
    endrule

    rule test_rule_376 (count >= 376);
        count <= count + 376;
        $display ("Executing Rule376");
    endrule

    rule test_rule_377 (count >= 377);
        count <= count + 377;
        $display ("Executing Rule377");
    endrule

    rule test_rule_378 (count >= 378);
        count <= count + 378;
        $display ("Executing Rule378");
    endrule

    rule test_rule_379 (count >= 379);
        count <= count + 379;
        $display ("Executing Rule379");
    endrule


    rule test_rule_380 (count >= 380);
        count <= count + 380;
        $display ("Executing Rule380");
    endrule

    rule test_rule_381 (count >= 381);
        count <= count + 381;
        $display ("Executing Rule381");
    endrule

    rule test_rule_382 (count >= 382);
        count <= count + 382;
        $display ("Executing Rule382");
    endrule

    rule test_rule_383 (count >= 383);
        count <= count + 383;
        $display ("Executing Rule383");
    endrule

    rule test_rule_384 (count >= 384);
        count <= count + 384;
        $display ("Executing Rule384");
    endrule

    rule test_rule_385 (count >= 385);
        count <= count + 385;
        $display ("Executing Rule385");
    endrule

    rule test_rule_386 (count >= 386);
        count <= count + 386;
        $display ("Executing Rule386");
    endrule

    rule test_rule_387 (count >= 387);
        count <= count + 387;
        $display ("Executing Rule387");
    endrule

    rule test_rule_388 (count >= 388);
        count <= count + 388;
        $display ("Executing Rule388");
    endrule

    rule test_rule_389 (count >= 389);
        count <= count + 389;
        $display ("Executing Rule389");
    endrule


    rule test_rule_390 (count >= 390);
        count <= count + 390;
        $display ("Executing Rule390");
    endrule

    rule test_rule_391 (count >= 391);
        count <= count + 391;
        $display ("Executing Rule391");
    endrule

    rule test_rule_392 (count >= 392);
        count <= count + 392;
        $display ("Executing Rule392");
    endrule

    rule test_rule_393 (count >= 393);
        count <= count + 393;
        $display ("Executing Rule393");
    endrule

    rule test_rule_394 (count >= 394);
        count <= count + 394;
        $display ("Executing Rule394");
    endrule

    rule test_rule_395 (count >= 395);
        count <= count + 395;
        $display ("Executing Rule395");
    endrule

    rule test_rule_396 (count >= 396);
        count <= count + 396;
        $display ("Executing Rule396");
    endrule

    rule test_rule_397 (count >= 397);
        count <= count + 397;
        $display ("Executing Rule397");
    endrule

    rule test_rule_398 (count >= 398);
        count <= count + 398;
        $display ("Executing Rule398");
    endrule

    rule test_rule_399 (count >= 399);
        count <= count + 399;
        $display ("Executing Rule399");
    endrule


    rule test_rule_400 (count >= 400);
        count <= count + 400;
        $display ("Executing Rule400");
    endrule

    rule test_rule_401 (count >= 401);
        count <= count + 401;
        $display ("Executing Rule401");
    endrule

    rule test_rule_402 (count >= 402);
        count <= count + 402;
        $display ("Executing Rule402");
    endrule

    rule test_rule_403 (count >= 403);
        count <= count + 403;
        $display ("Executing Rule403");
    endrule

    rule test_rule_404 (count >= 404);
        count <= count + 404;
        $display ("Executing Rule404");
    endrule

    rule test_rule_405 (count >= 405);
        count <= count + 405;
        $display ("Executing Rule405");
    endrule

    rule test_rule_406 (count >= 406);
        count <= count + 406;
        $display ("Executing Rule406");
    endrule

    rule test_rule_407 (count >= 407);
        count <= count + 407;
        $display ("Executing Rule407");
    endrule

    rule test_rule_408 (count >= 408);
        count <= count + 408;
        $display ("Executing Rule408");
    endrule

    rule test_rule_409 (count >= 409);
        count <= count + 409;
        $display ("Executing Rule409");
    endrule

    rule test_rule_410 (count >= 410);
        count <= count + 410;
        $display ("Executing Rule410");
    endrule

    rule test_rule_411 (count >= 411);
        count <= count + 411;
        $display ("Executing Rule411");
    endrule

    rule test_rule_412 (count >= 412);
        count <= count + 412;
        $display ("Executing Rule412");
    endrule

    rule test_rule_413 (count >= 413);
        count <= count + 413;
        $display ("Executing Rule413");
    endrule

    rule test_rule_414 (count >= 414);
        count <= count + 414;
        $display ("Executing Rule414");
    endrule

    rule test_rule_415 (count >= 415);
        count <= count + 415;
        $display ("Executing Rule415");
    endrule

    rule test_rule_416 (count >= 416);
        count <= count + 416;
        $display ("Executing Rule416");
    endrule

    rule test_rule_417 (count >= 417);
        count <= count + 417;
        $display ("Executing Rule417");
    endrule

    rule test_rule_418 (count >= 418);
        count <= count + 418;
        $display ("Executing Rule418");
    endrule

    rule test_rule_419 (count >= 419);
        count <= count + 419;
        $display ("Executing Rule419");
    endrule

    rule test_rule_420 (count >= 420);
        count <= count + 420;
        $display ("Executing Rule420");
    endrule

    rule test_rule_421 (count >= 421);
        count <= count + 421;
        $display ("Executing Rule421");
    endrule

    rule test_rule_422 (count >= 422);
        count <= count + 422;
        $display ("Executing Rule422");
    endrule

    rule test_rule_423 (count >= 423);
        count <= count + 423;
        $display ("Executing Rule423");
    endrule

    rule test_rule_424 (count >= 424);
        count <= count + 424;
        $display ("Executing Rule424");
    endrule

    rule test_rule_425 (count >= 425);
        count <= count + 425;
        $display ("Executing Rule425");
    endrule

    rule test_rule_426 (count >= 426);
        count <= count + 426;
        $display ("Executing Rule426");
    endrule

    rule test_rule_427 (count >= 427);
        count <= count + 427;
        $display ("Executing Rule427");
    endrule

    rule test_rule_428 (count >= 428);
        count <= count + 428;
        $display ("Executing Rule428");
    endrule

    rule test_rule_429 (count >= 429);
        count <= count + 429;
        $display ("Executing Rule429");
    endrule

    rule test_rule_430 (count >= 430);
        count <= count + 430;
        $display ("Executing Rule430");
    endrule

    rule test_rule_431 (count >= 431);
        count <= count + 431;
        $display ("Executing Rule431");
    endrule

    rule test_rule_432 (count >= 432);
        count <= count + 432;
        $display ("Executing Rule432");
    endrule

    rule test_rule_433 (count >= 433);
        count <= count + 433;
        $display ("Executing Rule433");
    endrule

    rule test_rule_434 (count >= 434);
        count <= count + 434;
        $display ("Executing Rule434");
    endrule

    rule test_rule_435 (count >= 435);
        count <= count + 435;
        $display ("Executing Rule435");
    endrule

    rule test_rule_436 (count >= 436);
        count <= count + 436;
        $display ("Executing Rule436");
    endrule

    rule test_rule_437 (count >= 437);
        count <= count + 437;
        $display ("Executing Rule437");
    endrule

    rule test_rule_438 (count >= 438);
        count <= count + 438;
        $display ("Executing Rule438");
    endrule

    rule test_rule_439 (count >= 439);
        count <= count + 439;
        $display ("Executing Rule439");
    endrule


    rule test_rule_440 (count >= 440);
        count <= count + 440;
        $display ("Executing Rule440");
    endrule

    rule test_rule_441 (count >= 441);
        count <= count + 441;
        $display ("Executing Rule441");
    endrule

    rule test_rule_442 (count >= 442);
        count <= count + 442;
        $display ("Executing Rule442");
    endrule

    rule test_rule_443 (count >= 443);
        count <= count + 443;
        $display ("Executing Rule443");
    endrule

    rule test_rule_444 (count >= 444);
        count <= count + 444;
        $display ("Executing Rule444");
    endrule

    rule test_rule_445 (count >= 445);
        count <= count + 445;
        $display ("Executing Rule445");
    endrule

    rule test_rule_446 (count >= 446);
        count <= count + 446;
        $display ("Executing Rule446");
    endrule

    rule test_rule_447 (count >= 447);
        count <= count + 447;
        $display ("Executing Rule447");
    endrule

    rule test_rule_448 (count >= 448);
        count <= count + 448;
        $display ("Executing Rule448");
    endrule

    rule test_rule_449 (count >= 449);
        count <= count + 449;
        $display ("Executing Rule449");
    endrule


    rule test_rule_450 (count >= 450);
        count <= count + 450;
        $display ("Executing Rule450");
    endrule

    rule test_rule_451 (count >= 451);
        count <= count + 451;
        $display ("Executing Rule451");
    endrule

    rule test_rule_452 (count >= 452);
        count <= count + 452;
        $display ("Executing Rule452");
    endrule

    rule test_rule_453 (count >= 453);
        count <= count + 453;
        $display ("Executing Rule453");
    endrule

    rule test_rule_454 (count >= 454);
        count <= count + 454;
        $display ("Executing Rule454");
    endrule

    rule test_rule_455 (count >= 455);
        count <= count + 455;
        $display ("Executing Rule455");
    endrule

    rule test_rule_456 (count >= 456);
        count <= count + 456;
        $display ("Executing Rule456");
    endrule

    rule test_rule_457 (count >= 457);
        count <= count + 457;
        $display ("Executing Rule457");
    endrule

    rule test_rule_458 (count >= 458);
        count <= count + 458;
        $display ("Executing Rule458");
    endrule

    rule test_rule_459 (count >= 459);
        count <= count + 459;
        $display ("Executing Rule459");
    endrule


    rule test_rule_460 (count >= 460);
        count <= count + 460;
        $display ("Executing Rule460");
    endrule

    rule test_rule_461 (count >= 461);
        count <= count + 461;
        $display ("Executing Rule461");
    endrule

    rule test_rule_462 (count >= 462);
        count <= count + 462;
        $display ("Executing Rule462");
    endrule

    rule test_rule_463 (count >= 463);
        count <= count + 463;
        $display ("Executing Rule463");
    endrule

    rule test_rule_464 (count >= 464);
        count <= count + 464;
        $display ("Executing Rule464");
    endrule

    rule test_rule_465 (count >= 465);
        count <= count + 465;
        $display ("Executing Rule465");
    endrule

    rule test_rule_466 (count >= 466);
        count <= count + 466;
        $display ("Executing Rule466");
    endrule

    rule test_rule_467 (count >= 467);
        count <= count + 467;
        $display ("Executing Rule467");
    endrule

    rule test_rule_468 (count >= 468);
        count <= count + 468;
        $display ("Executing Rule468");
    endrule

    rule test_rule_469 (count >= 469);
        count <= count + 469;
        $display ("Executing Rule469");
    endrule


    rule test_rule_470 (count >= 470);
        count <= count + 470;
        $display ("Executing Rule470");
    endrule

    rule test_rule_471 (count >= 471);
        count <= count + 471;
        $display ("Executing Rule471");
    endrule

    rule test_rule_472 (count >= 472);
        count <= count + 472;
        $display ("Executing Rule472");
    endrule

    rule test_rule_473 (count >= 473);
        count <= count + 473;
        $display ("Executing Rule473");
    endrule

    rule test_rule_474 (count >= 474);
        count <= count + 474;
        $display ("Executing Rule474");
    endrule

    rule test_rule_475 (count >= 475);
        count <= count + 475;
        $display ("Executing Rule475");
    endrule

    rule test_rule_476 (count >= 476);
        count <= count + 476;
        $display ("Executing Rule476");
    endrule

    rule test_rule_477 (count >= 477);
        count <= count + 477;
        $display ("Executing Rule477");
    endrule

    rule test_rule_478 (count >= 478);
        count <= count + 478;
        $display ("Executing Rule478");
    endrule

    rule test_rule_479 (count >= 479);
        count <= count + 479;
        $display ("Executing Rule479");
    endrule


    rule test_rule_480 (count >= 480);
        count <= count + 480;
        $display ("Executing Rule480");
    endrule

    rule test_rule_481 (count >= 481);
        count <= count + 481;
        $display ("Executing Rule481");
    endrule

    rule test_rule_482 (count >= 482);
        count <= count + 482;
        $display ("Executing Rule482");
    endrule

    rule test_rule_483 (count >= 483);
        count <= count + 483;
        $display ("Executing Rule483");
    endrule

    rule test_rule_484 (count >= 484);
        count <= count + 484;
        $display ("Executing Rule484");
    endrule

    rule test_rule_485 (count >= 485);
        count <= count + 485;
        $display ("Executing Rule485");
    endrule

    rule test_rule_486 (count >= 486);
        count <= count + 486;
        $display ("Executing Rule486");
    endrule

    rule test_rule_487 (count >= 487);
        count <= count + 487;
        $display ("Executing Rule487");
    endrule

    rule test_rule_488 (count >= 488);
        count <= count + 488;
        $display ("Executing Rule488");
    endrule

    rule test_rule_489 (count >= 489);
        count <= count + 489;
        $display ("Executing Rule489");
    endrule


    rule test_rule_490 (count >= 490);
        count <= count + 490;
        $display ("Executing Rule490");
    endrule

    rule test_rule_491 (count >= 491);
        count <= count + 491;
        $display ("Executing Rule491");
    endrule

    rule test_rule_492 (count >= 492);
        count <= count + 492;
        $display ("Executing Rule492");
    endrule

    rule test_rule_493 (count >= 493);
        count <= count + 493;
        $display ("Executing Rule493");
    endrule

    rule test_rule_494 (count >= 494);
        count <= count + 494;
        $display ("Executing Rule494");
    endrule

    rule test_rule_495 (count >= 495);
        count <= count + 495;
        $display ("Executing Rule495");
    endrule

    rule test_rule_496 (count >= 496);
        count <= count + 496;
        $display ("Executing Rule496");
    endrule

    rule test_rule_497 (count >= 497);
        count <= count + 497;
        $display ("Executing Rule497");
    endrule

    rule test_rule_498 (count >= 498);
        count <= count + 498;
        $display ("Executing Rule498");
    endrule

    rule test_rule_499 (count >= 499);
        count <= count + 499;
        $display ("Executing Rule499");
    endrule

    rule test_rule_500 (count >= 500);
        count <= count + 500;
        $display ("Executing Rule500");
    endrule








    rule always_schedule (True);
         count2 <= count2 + 1;
    endrule

    rule endsim (count2 == 2047);
        $finish (2'b00);
    endrule

endmodule : mkFive_Hundred_Rules

endpackage : Five_Hundred_Rules
