Bit #(10) tenBits;
tenBits = 10;

Bit #(2) twoBits;
twoBits = tenBits[1:0];

Bit #(3) threeBits;
threeBits = tenBits[8:6];
