typeclass Foo#(type x)
 dependencies (x determines y);
   function y fooFn(x x1);
endtypeclass
