interface Test;
 method Bit#(1) out(Bit#(1) in);
endinterface: Test
