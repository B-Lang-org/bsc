function int f(Bool x);
   (* foo *)
   case (x)
      True: return 1;
      False: return 2;
   endcase
endfunction

