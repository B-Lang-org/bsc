package NumWhereNonNumExpected () where

data (Foo :: * -> *) a = Bar a

x :: Foo 1
x = 0

