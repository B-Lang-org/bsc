module mkProvisoProvisoMismatch_TopLevel(Reg#(t))
   provisos(Bits#(szt, j), Bits#(t, szt));
endmodule
