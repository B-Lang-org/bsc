import FIFO :: * ;
import FIFOLevel :: *;

`include "FIFO.include.bsv"
`include "FIFOLevel.include.bsv"

