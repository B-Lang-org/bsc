-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EBadModuleInterface1.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers a "multiple interface expressions" error (EBadModuleInterface)

-- Error Message : bsc EBadModuleInterface1.bs
-- bsc: Compilation errors:
-- "EBadModuleInterface1.bs", line 26, column 4, Multiple interface expressions
-----------------------------------------------------------------------

package EBadModuleInterface1 (EBadModuleInterface1(..), mkEBadModuleInterface1) where

-- import Int

interface EBadModuleInterface1 =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32


mkEBadModuleInterface1 :: Module EBadModuleInterface1
mkEBadModuleInterface1 =
    module

        x :: Reg (Int 32)
        x <- mkReg 0

	y :: Reg (Int 32)
	y <- mkReg 0

        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0


        interface
            start ix iy = action
                              x := ix
                              y := iy
                          when y == 0
            result = x when y == 0

