package StmtBind_NoType () where

x :: Module Empty
x = module
      _ <- mkReg True

      interface {}

