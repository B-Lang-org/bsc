package TestCShow where

import CShow
import ListN
import Vector
import BuildVector

data Foo = A (UInt 8) Bool Bar
         | B (Int 16)
         | C
         | D {a :: (Bit 8); b :: Foo}
  deriving (FShow)

struct Bar =
  foo :: Foo
  x :: (UInt 8)
 deriving (FShow)

data Baz a = Baz a a
  deriving (FShow)

sysTestCShow :: Module Empty
sysTestCShow = module
  rules
    when True ==> do
      $display (cshow (42 :: UInt 8))
      $display (cshow (3.14 :: Real))
      $display (cshow '*')
      $display (cshow "Hello")
      $display (cshow $ $format "Hello")
      $display (cshow ())
      $display (cshow (Bar {x=42; foo=C}))
      $display (cshow (A 12 True (Bar {foo=D {a=34; b=C}; x=42})))
      $display (cshow (Baz C (A 12 True (Bar {foo=D {a=34; b=C}; x=42}))))
      $display (cshow ((vec (Bar {x=42; foo=C}) (Bar {x=3; foo=B 2323})) :: Vector 2 Bar))
      $display (cshow ((Bar {x=42; foo=C}) :> (Bar {x=3; foo=B 2323}) :> ListN.nil))
      $display (cshow ("x", ((Left 123) :: Either (UInt 8) Bar, False)))
      $finish
