package Math;

import Complex::*;
import FixedPoint::*;
import NumberTypes::*;
import Divide::*;
import SquareRoot::*;
import FloatingPoint::*;

endpackage
