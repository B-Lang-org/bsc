package EWeakContext2() where

foo :: a
foo = 0

