/*
PURPOSE - Simple testcase using the 'define preprocessor directive
 
*/
package Design ;

import Vector::*;



function Bit#(4) result (Bit #(4) x);
`define max 23
Bit #(4) res;
  res = x ^ (x >> 1) ;
  return res;
endfunction 


endpackage