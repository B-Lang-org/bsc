package PackageEmpty;
endpackage: PackageEmpty
