package StmtBind_Type_OneLine () where

x :: Module Empty
x = module
      _ :: Reg Bool <- mkReg True

      interface {}

