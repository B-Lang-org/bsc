`define is 1
`define fs 5
`define full sysFromReal_1_5

`include "FromReal.bsv"
