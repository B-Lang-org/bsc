package FShow;

// The FShow typeclass is now defined in the Prelude and FShow instances
// are defined alongside the types, so there is no need for this file.
// However, we provide this empty package, so that existing code that
// imports the FShow package will still compile.

endpackage

