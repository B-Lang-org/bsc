-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EUnboundTyCon.bs

-- Author : Nitin Chand Rahul <ncr@noida.interrasystems.com>

-- Description: This testcase triggers the EUnboundTyCon error of the bluespec
-- compiler (Unbound Type Constructor)
--
-----------------------------------------------------------------------



package EUnboundTyCon () where

interface GCD =
    start  :: R 32 -> R 32 -> Action  -- Type Constructor R not bounded
    result :: R 32

mkGCD :: Module GCD
mkGCD =
    module
	x :: Reg (R 32)
	x <- mkRegU

	y :: Reg (R 32)
	y <- mkReg 0

        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0


