(* synthesize *)
module sysPrintType3();

  messageM(printType(typeOf(Nothing)));

endmodule

