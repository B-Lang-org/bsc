package LevelFIFO ;

import FIFOLevel:: *;

export FIFOLevel :: *;


endpackage
