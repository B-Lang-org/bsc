function bit[3:0] f();
  return 3;
endfunction
