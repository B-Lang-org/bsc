import Vector::*;

(* synthesize *)
module sysInvalidPortName ( (* port="hey mom!" *)Vector#(2,Bool) xs,
                            Empty ifc);
endmodule

