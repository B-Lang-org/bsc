typeclass C #(type a, type b, type a);
  function Action fn(a v1, b v2);
endtypeclass
