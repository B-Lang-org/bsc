
(* always_ready = "foo,bar,Bat" *)
module sysT2();
endmodule

