(* synthesize *)
module sysShowVersionTimestamps ();
  rule r;
    $display("Success");
    $finish(0);
  endrule
endmodule

