(* synthesize *)
(* default_clock_osc = "clk" *)
module sysRenamedClockClash();
endmodule
