`define foo // This is a commment \