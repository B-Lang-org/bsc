(* synthesize *)
module sysOctalCharsAsInteger();
rule test;
$display(primStringToInteger("\000"));
$display(primStringToInteger("\001"));
$display(primStringToInteger("\002"));
$display(primStringToInteger("\003"));
$display(primStringToInteger("\004"));
$display(primStringToInteger("\005"));
$display(primStringToInteger("\006"));
$display(primStringToInteger("\007"));
$display(primStringToInteger("\010"));
$display(primStringToInteger("\011"));
$display(primStringToInteger("\012"));
$display(primStringToInteger("\013"));
$display(primStringToInteger("\014"));
$display(primStringToInteger("\015"));
$display(primStringToInteger("\016"));
$display(primStringToInteger("\017"));
$display(primStringToInteger("\020"));
$display(primStringToInteger("\021"));
$display(primStringToInteger("\022"));
$display(primStringToInteger("\023"));
$display(primStringToInteger("\024"));
$display(primStringToInteger("\025"));
$display(primStringToInteger("\026"));
$display(primStringToInteger("\027"));
$display(primStringToInteger("\030"));
$display(primStringToInteger("\031"));
$display(primStringToInteger("\032"));
$display(primStringToInteger("\033"));
$display(primStringToInteger("\034"));
$display(primStringToInteger("\035"));
$display(primStringToInteger("\036"));
$display(primStringToInteger("\037"));
$display(primStringToInteger("\040"));
$display(primStringToInteger("\041"));
$display(primStringToInteger("\042"));
$display(primStringToInteger("\043"));
$display(primStringToInteger("\044"));
$display(primStringToInteger("\045"));
$display(primStringToInteger("\046"));
$display(primStringToInteger("\047"));
$display(primStringToInteger("\050"));
$display(primStringToInteger("\051"));
$display(primStringToInteger("\052"));
$display(primStringToInteger("\053"));
$display(primStringToInteger("\054"));
$display(primStringToInteger("\055"));
$display(primStringToInteger("\056"));
$display(primStringToInteger("\057"));
$display(primStringToInteger("\060"));
$display(primStringToInteger("\061"));
$display(primStringToInteger("\062"));
$display(primStringToInteger("\063"));
$display(primStringToInteger("\064"));
$display(primStringToInteger("\065"));
$display(primStringToInteger("\066"));
$display(primStringToInteger("\067"));
$display(primStringToInteger("\070"));
$display(primStringToInteger("\071"));
$display(primStringToInteger("\072"));
$display(primStringToInteger("\073"));
$display(primStringToInteger("\074"));
$display(primStringToInteger("\075"));
$display(primStringToInteger("\076"));
$display(primStringToInteger("\077"));
$display(primStringToInteger("\100"));
$display(primStringToInteger("\101"));
$display(primStringToInteger("\102"));
$display(primStringToInteger("\103"));
$display(primStringToInteger("\104"));
$display(primStringToInteger("\105"));
$display(primStringToInteger("\106"));
$display(primStringToInteger("\107"));
$display(primStringToInteger("\110"));
$display(primStringToInteger("\111"));
$display(primStringToInteger("\112"));
$display(primStringToInteger("\113"));
$display(primStringToInteger("\114"));
$display(primStringToInteger("\115"));
$display(primStringToInteger("\116"));
$display(primStringToInteger("\117"));
$display(primStringToInteger("\120"));
$display(primStringToInteger("\121"));
$display(primStringToInteger("\122"));
$display(primStringToInteger("\123"));
$display(primStringToInteger("\124"));
$display(primStringToInteger("\125"));
$display(primStringToInteger("\126"));
$display(primStringToInteger("\127"));
$display(primStringToInteger("\130"));
$display(primStringToInteger("\131"));
$display(primStringToInteger("\132"));
$display(primStringToInteger("\133"));
$display(primStringToInteger("\134"));
$display(primStringToInteger("\135"));
$display(primStringToInteger("\136"));
$display(primStringToInteger("\137"));
$display(primStringToInteger("\140"));
$display(primStringToInteger("\141"));
$display(primStringToInteger("\142"));
$display(primStringToInteger("\143"));
$display(primStringToInteger("\144"));
$display(primStringToInteger("\145"));
$display(primStringToInteger("\146"));
$display(primStringToInteger("\147"));
$display(primStringToInteger("\150"));
$display(primStringToInteger("\151"));
$display(primStringToInteger("\152"));
$display(primStringToInteger("\153"));
$display(primStringToInteger("\154"));
$display(primStringToInteger("\155"));
$display(primStringToInteger("\156"));
$display(primStringToInteger("\157"));
$display(primStringToInteger("\160"));
$display(primStringToInteger("\161"));
$display(primStringToInteger("\162"));
$display(primStringToInteger("\163"));
$display(primStringToInteger("\164"));
$display(primStringToInteger("\165"));
$display(primStringToInteger("\166"));
$display(primStringToInteger("\167"));
$display(primStringToInteger("\170"));
$display(primStringToInteger("\171"));
$display(primStringToInteger("\172"));
$display(primStringToInteger("\173"));
$display(primStringToInteger("\174"));
$display(primStringToInteger("\175"));
$display(primStringToInteger("\176"));
$display(primStringToInteger("\177"));
$display(primStringToInteger("\200"));
$display(primStringToInteger("\201"));
$display(primStringToInteger("\202"));
$display(primStringToInteger("\203"));
$display(primStringToInteger("\204"));
$display(primStringToInteger("\205"));
$display(primStringToInteger("\206"));
$display(primStringToInteger("\207"));
$display(primStringToInteger("\210"));
$display(primStringToInteger("\211"));
$display(primStringToInteger("\212"));
$display(primStringToInteger("\213"));
$display(primStringToInteger("\214"));
$display(primStringToInteger("\215"));
$display(primStringToInteger("\216"));
$display(primStringToInteger("\217"));
$display(primStringToInteger("\220"));
$display(primStringToInteger("\221"));
$display(primStringToInteger("\222"));
$display(primStringToInteger("\223"));
$display(primStringToInteger("\224"));
$display(primStringToInteger("\225"));
$display(primStringToInteger("\226"));
$display(primStringToInteger("\227"));
$display(primStringToInteger("\230"));
$display(primStringToInteger("\231"));
$display(primStringToInteger("\232"));
$display(primStringToInteger("\233"));
$display(primStringToInteger("\234"));
$display(primStringToInteger("\235"));
$display(primStringToInteger("\236"));
$display(primStringToInteger("\237"));
$display(primStringToInteger("\240"));
$display(primStringToInteger("\241"));
$display(primStringToInteger("\242"));
$display(primStringToInteger("\243"));
$display(primStringToInteger("\244"));
$display(primStringToInteger("\245"));
$display(primStringToInteger("\246"));
$display(primStringToInteger("\247"));
$display(primStringToInteger("\250"));
$display(primStringToInteger("\251"));
$display(primStringToInteger("\252"));
$display(primStringToInteger("\253"));
$display(primStringToInteger("\254"));
$display(primStringToInteger("\255"));
$display(primStringToInteger("\256"));
$display(primStringToInteger("\257"));
$display(primStringToInteger("\260"));
$display(primStringToInteger("\261"));
$display(primStringToInteger("\262"));
$display(primStringToInteger("\263"));
$display(primStringToInteger("\264"));
$display(primStringToInteger("\265"));
$display(primStringToInteger("\266"));
$display(primStringToInteger("\267"));
$display(primStringToInteger("\270"));
$display(primStringToInteger("\271"));
$display(primStringToInteger("\272"));
$display(primStringToInteger("\273"));
$display(primStringToInteger("\274"));
$display(primStringToInteger("\275"));
$display(primStringToInteger("\276"));
$display(primStringToInteger("\277"));
$display(primStringToInteger("\300"));
$display(primStringToInteger("\301"));
$display(primStringToInteger("\302"));
$display(primStringToInteger("\303"));
$display(primStringToInteger("\304"));
$display(primStringToInteger("\305"));
$display(primStringToInteger("\306"));
$display(primStringToInteger("\307"));
$display(primStringToInteger("\310"));
$display(primStringToInteger("\311"));
$display(primStringToInteger("\312"));
$display(primStringToInteger("\313"));
$display(primStringToInteger("\314"));
$display(primStringToInteger("\315"));
$display(primStringToInteger("\316"));
$display(primStringToInteger("\317"));
$display(primStringToInteger("\320"));
$display(primStringToInteger("\321"));
$display(primStringToInteger("\322"));
$display(primStringToInteger("\323"));
$display(primStringToInteger("\324"));
$display(primStringToInteger("\325"));
$display(primStringToInteger("\326"));
$display(primStringToInteger("\327"));
$display(primStringToInteger("\330"));
$display(primStringToInteger("\331"));
$display(primStringToInteger("\332"));
$display(primStringToInteger("\333"));
$display(primStringToInteger("\334"));
$display(primStringToInteger("\335"));
$display(primStringToInteger("\336"));
$display(primStringToInteger("\337"));
$display(primStringToInteger("\340"));
$display(primStringToInteger("\341"));
$display(primStringToInteger("\342"));
$display(primStringToInteger("\343"));
$display(primStringToInteger("\344"));
$display(primStringToInteger("\345"));
$display(primStringToInteger("\346"));
$display(primStringToInteger("\347"));
$display(primStringToInteger("\350"));
$display(primStringToInteger("\351"));
$display(primStringToInteger("\352"));
$display(primStringToInteger("\353"));
$display(primStringToInteger("\354"));
$display(primStringToInteger("\355"));
$display(primStringToInteger("\356"));
$display(primStringToInteger("\357"));
$display(primStringToInteger("\360"));
$display(primStringToInteger("\361"));
$display(primStringToInteger("\362"));
$display(primStringToInteger("\363"));
$display(primStringToInteger("\364"));
$display(primStringToInteger("\365"));
$display(primStringToInteger("\366"));
$display(primStringToInteger("\367"));
$display(primStringToInteger("\370"));
$display(primStringToInteger("\371"));
$display(primStringToInteger("\372"));
$display(primStringToInteger("\373"));
$display(primStringToInteger("\374"));
$display(primStringToInteger("\375"));
$display(primStringToInteger("\376"));
$display(primStringToInteger("\377"));
$finish(0);
endrule
endmodule
