import Vector::*;

(* synthesize *)
(* gate_all_clocks *)
module sysGateAllClocks_VecClock ( Vector#(2,Clock) clks,
                                   Empty ifc );
endmodule

