function Bool f(a#(4) y);
  a#(Bool) x = ?;
  return True;
endfunction


