
(* always_ready = "start" *)
interface Ifc;
  method Action start(Bool a, Bool b);
endinterface

