let _ = True;
