
export x;
export x;
export x;

Bool x = True;

