package TypeAliasParamGivenTooMany_OK () where

type (Foo :: # -> *) = Bit

