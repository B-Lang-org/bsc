(* synthesize *)
module sysDontCareFmt();

   rule rl;
      Fmt f = ?;
      $display(f);
   endrule

endmodule

