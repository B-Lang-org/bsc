package DataDefFieldIsNum () where

data Foo = Bar 12

