-----------------------------------------------------------------------
-- Project: Bluespec

-- File: ERTSHeapExhausted1.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers a "Out of Heap" error by the Run Time System
-- For the current test-case this message will be generated for all selections of
-- maximum Heap less than 1 MB  Ex.. M256k , M512k etc.

-- Error Message : bsc +RTS -M1M -RTS -verilog -g mkERTSHeapExhausted1 ERTSHeapExhausted1.bs
-- Heap exhausted;
-- Current maximum heap size is 999424 bytes;
-- use `+RTS -M<size>' to increase it.

-----------------------------------------------------------------------

package ERTSHeapExhausted1 (ERTSHeapExhausted1(..), mkERTSHeapExhausted1) where

-- import Int

interface ERTSHeapExhausted1 =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32

mkERTSHeapExhausted1 :: Module ERTSHeapExhausted1
mkERTSHeapExhausted1 =
    module
	x :: Reg (Int 32)
	x <- mkRegU

	y :: Reg (Int 32)
	y <- mkReg 0

        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0


