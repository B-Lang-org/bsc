package ReExportSame_Top;

import ReExportSame_P::*;
import ReExportSame_Sub::*;

export ReExportSame_P::*;
export ReExportSame_Sub::*;

endpackage

