function Action f();
  action
    return ?;
  endaction
endfunction
