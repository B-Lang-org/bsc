typedef enum { A, B }
  AB deriving(Eq,Bits);

AB a = A;

AB b = B;

