
interface Ifc;
 (* result = "always" *)
 method Bool check ();
endinterface

(* synthesize *)
module mkKeyword (Ifc);
endmodule
