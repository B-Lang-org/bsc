package ExclusiveEnq (sysExclusiveEnq) where

import FIFO

sysExclusiveEnq :: Module Empty
sysExclusiveEnq =
  module
    f :: FIFO (Bit 3) <- mkFIFO
    b :: Reg (Bool)  <- mkReg False
    counter :: Reg (Bit 5) <- mkReg 0

    rules
      when True ==>
         b := not b
      when True ==>
         action
           if b then f.enq 5 else noAction
           if not b then f.enq 7 else noAction
      when True ==>
         if (counter > 10) then $finish 0 else $display "%0d" (1 :: Bit 3)
      when True ==> counter := counter + 1

