package TypeAliasResGivenNumIsNonNum () where

type (Foo :: # -> #) a = Bit a

