package NoSign where

x = 17
