package TwoArgMissingOne () where

data Foo a b = Bar a b

x :: Foo Bool
x = _

