function Bool f();
  int y;
  for (int x=1, y=0, int z=3; x<3; x=x+1)
  begin
    y = y + x;
  end
  return False;
endfunction
