package ReExportSame_TopBad2;

import ReExportSame_P::*;
import ReExportSame_Q::*;

export ReExportSame_P::*;
export ReExportSame_Q::*;

endpackage

