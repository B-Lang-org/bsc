function bit[3:0] f(Bool cond);
  if (cond)
    return 3;
  else
    return 5;
endfunction
