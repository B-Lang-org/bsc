module sysAmbigTCon_TLog (Reg#(Bit#(TLog#(n))));
endmodule
