Bit#(8) x = truncate(1);
