function Action f();
   action
      (* foo *)
      noAction;
   endaction
endfunction

