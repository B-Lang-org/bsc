
function a#(m) x(a#(m) y) provisos (BitExtend#(n,m,a));
   return (truncate(zeroExtend(y)));
endfunction

