package ExportAllImportBad where

import ExportAllExportBad

quux :: Bool
quux = foo || bar
