module mkFoo();
  Reg#(Bool) r <- mkRegU();
endmodule
