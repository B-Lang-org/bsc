typedef union tagged { Bool Foo; } Bar;

Bar x = Foo;

