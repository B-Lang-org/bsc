package ShallowSplit where

import Vector
import BuildVector
import SplitPorts
import CShow

struct Foo =
  x :: Int 8
  y :: Int 8
 deriving (Bits)

struct Bar =
  v :: Vector 3 Bool
  w :: (Bool, UInt 16)
  z :: Foo
 deriving (Bits)

struct Baz =
  a :: Maybe Foo
  b :: Bar
  c :: Vector 3 (Vector 8 Foo, Bar)
  d :: ()
  e :: Vector 0 Foo
 -- No Bits instance needed

interface SplitTest =
  putFoo :: ShallowSplit Foo -> Action
  putBar :: ShallowSplit Bar -> Action {-# prefix = "PUT_BAR" #-}
  putFooBar :: ShallowSplit Foo -> ShallowSplit Bar -> Action {-# arg_names = ["fooIn", "barIn"] #-}
  putFoos :: ShallowSplit (Vector 50 Foo) -> Action
  putBaz :: ShallowSplit Baz -> Action

  getFoo :: ShallowSplit Foo
  getBar :: ShallowSplit Foo -> ShallowSplit Bar {-# result = "GET_BAR" #-}

  update :: ShallowSplit Foo -> ActionValue (ShallowSplit Bar)


{-# synthesize mkShallowSplitTest #-}
mkShallowSplitTest :: Module SplitTest
mkShallowSplitTest =
  module
    theCond <- mkReg False
    theFoo <- mkReg (Foo { x = 0; y = 0; })
    interface
      putFoo (ShallowSplit x) = $display "putFoo: " (cshow x)
      putBar (ShallowSplit x) = $display "putBar: " (cshow x)
      putFooBar (ShallowSplit x) (ShallowSplit y) = $display "putFooBar: " (cshow x) " " (cshow y)
      putFoos (ShallowSplit x) = $display "putFoos: " (cshow x)
      putBaz (ShallowSplit x) = $display "putBaz: " (cshow x)
      getFoo = ShallowSplit $ Foo { x = 42; y = 43; }
      getBar (ShallowSplit f) = ShallowSplit $ Bar { v = vec True False True; w = (False, 0x4321); z = f; }
      update (ShallowSplit f) = do
        theCond := not theCond
        theFoo := f
        return $ ShallowSplit $ Bar { v = vec (f.x == 33) theCond (not theCond); w = (theCond, 0xDEAD); z = theFoo; }

{-# synthesize sysShallowSplit #-}
sysShallowSplit :: Module Empty
sysShallowSplit =
  module
    s <- mkShallowSplitTest
    i :: Reg (UInt 8) <- mkReg 0
    rules
      when True ==> i := i + 1
      when i == 0 ==> s.putFoo $ ShallowSplit $ Foo { x = 1; y = 2; }
      when i == 1 ==> s.putBar $ ShallowSplit $ Bar { v = vec True False True; w = (True, 0x1234); z = Foo { x = 3; y = 4; } }
      when i == 2 ==> s.putFooBar (ShallowSplit $ Foo { x = 5; y = 6; }) (ShallowSplit $ Bar { v = vec False True False; w = (False, 0x5678); z = Foo { x = 7; y = 8; } })
      when i == 3 ==> s.putFoos $ ShallowSplit $ genWith $ \ j -> Foo { x = fromInteger $ 9 + j / 2; y = fromInteger $ 10 - 2*j / 3; }
      when i == 4 ==> s.putBaz $ ShallowSplit $ Baz { a = Just $ Foo { x = 9; y = 10; }; b = Bar { v = vec True False False; w = (True, 0x1234); z = Foo { x = 3; y = 4; }; }; c = vec (vec (Foo { x = 11; y = 12; }) (Foo { x = 13; y = 14; }) (Foo { x = 15; y = 16; }) (Foo { x = 17; y = 18; }) (Foo { x = 19; y = 20; }) (Foo { x = 21; y = 22; }) (Foo { x = 23; y = 24; }) (Foo { x = 25; y = 26; }), Bar { v = vec True False True; w = (True, 0xBEEF); z = Foo { x = 3; y = 4; } }) (vec (Foo { x = 27; y = 28; }) (Foo { x = 29; y = 30; }) (Foo { x = 31; y = 32; }) (Foo { x = 33; y = 34; }) (Foo { x = 35; y = 36; }) (Foo { x = 37; y = 38; }) (Foo { x = 39; y = 40; }) (Foo { x = 41; y = 42; }), Bar { v = vec True False True; w = (True, 0x4321); z = Foo { x = 123; y = 42; } }) (vec (Foo { x = 43; y = 44; }) (Foo { x = 45; y = 46; }) (Foo { x = 47; y = 48; }) (Foo { x = 49; y = 50; }) (Foo { x = 51; y = 52; }) (Foo { x = 53; y = 54; }) (Foo { x = 55; y = 56; }) (Foo { x = 57; y = 58; }), Bar { v = vec True True True; w = (True, 0xAABB); z = Foo { x = 3; y = 4; } }); d = (); e = nil; }
      when i == 5 ==> $display "getFoo: " (cshow s.getFoo)
      when i == 6 ==> $display "getBar: " (cshow $ s.getBar s.getFoo)
      when i == 7 ==> do
        res <- s.update (ShallowSplit $ Foo { x = 77; y = 88; })
        $display "update: " (cshow res)
      when i == 8 ==> do
        res <- s.update (ShallowSplit $ Foo { x = 33; y = 44; })
        $display "update: " (cshow res)
      when i == 9 ==> $finish
