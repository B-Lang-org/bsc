-- Tests to explore the compiler's output for derived Bits instances.
package Alt5 where

data Alt5
    = A (Bit 1)
    | B
    | C (Bit 1)
    | D
    deriving (Bits)

interface TestTags =
  isA :: Bool
  isB :: Bool
  isC :: Bool
  isD :: Bool

{-# verilog mkAlt5Reg #-}
mkAlt5Reg :: Module (Reg Alt5)
mkAlt5Reg =
  module
    r <- mkRegU
    return r

{-# verilog mkMaybeAlt5Reg #-}
mkMaybeAlt5Reg :: Module (Reg (Maybe Alt5))
mkMaybeAlt5Reg =
  module
    r <- mkRegU
    return r

{-# verilog mkAlt5Test #-}
mkAlt5Test :: Module TestTags
mkAlt5Test =
  module
   r :: Reg Alt5 <- mkRegU
   interface TestTags
     isA = case r of
            A _ -> True
            _   -> False
     isB = case r of
            B   -> True
            _   -> False
     isC = case r of
            C _ -> True
            _   -> False
     isD = case r of
            D   -> True
            _   -> False
