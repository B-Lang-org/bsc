typedef Foo Bar;
typedef Bar Foo;

Foo x = 0;



