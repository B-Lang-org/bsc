package StringKindPolyToSpecific where

data (Foo :: $ -> *) s = Foo

a :: Foo a
a = Foo

b :: Foo "b"
b = a

