module sysAmbigTCon_TMul (Reg#(Bit#(TMul#(x,y))));
endmodule
