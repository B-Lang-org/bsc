function Bool fn(Bool _);
  return _;
endfunction
