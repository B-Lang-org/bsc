`define is 5
`define fs 1
`define full sysFromReal_5_1

`include "FromReal.bsv"
