package IfReadBug(sysIfReadBug) where

interface Foo a =
  read :: a -> a

{-# verilog mkFoo #-}
mkFoo :: Module (Foo (Bit 16))
mkFoo =
 module
   interface
     read x = x

sysIfReadBug :: Module Empty
sysIfReadBug =
  module
    r :: Reg (Bit 16) <- mkRegU
    f :: Foo (Bit 16) <- mkFoo
    b :: Reg (Bool) <- mkRegU

    rules
      when (True) ==>
       if b then
        r := f.read (0x0019)
       else
        r := f.read (0x0023)


