function int foo (int x) ;
        (* split *)
        if (x==10)
        return 20;
        else
        return 30;
endfunction
