interface Null;
endinterface

module mkEmpty(Null);
endmodule
