import RegFile::*;

interface InvSboxRom;
   method Bit#(8) read( Bit#(8) addr );
endinterface

(* synthesize, always_ready, always_enabled *)
module mkInvSboxRom ( InvSboxRom );
   method Bit#(8) read( Bit#(8) addr ) =
      case (addr)
         0: return 8'h52;
         1: return 8'h09;
         2: return 8'h6a;
         3: return 8'hd5;
         4: return 8'h30;
         5: return 8'h36;
         6: return 8'ha5;
         7: return 8'h38;
         8: return 8'hbf;
         9: return 8'h40;
         10: return 8'ha3;
         11: return 8'h9e;
         12: return 8'h81;
         13: return 8'hf3;
         14: return 8'hd7;
         15: return 8'hfb;
         16: return 8'h7c;
         17: return 8'he3;
         18: return 8'h39;
         19: return 8'h82;
         20: return 8'h9b;
         21: return 8'h2f;
         22: return 8'hff;
         23: return 8'h87;
         24: return 8'h34;
         25: return 8'h8e;
         26: return 8'h43;
         27: return 8'h44;
         28: return 8'hc4;
         29: return 8'hde;
         30: return 8'he9;
         31: return 8'hcb;
         32: return 8'h54;
         33: return 8'h7b;
         34: return 8'h94;
         35: return 8'h32;
         36: return 8'ha6;
         37: return 8'hc2;
         38: return 8'h23;
         39: return 8'h3d;
         40: return 8'hee;
         41: return 8'h4c;
         42: return 8'h95;
         43: return 8'h0b;
         44: return 8'h42;
         45: return 8'hfa;
         46: return 8'hc3;
         47: return 8'h4e;
         48: return 8'h08;
         49: return 8'h2e;
         50: return 8'ha1;
         51: return 8'h66;
         52: return 8'h28;
         53: return 8'hd9;
         54: return 8'h24;
         55: return 8'hb2;
         56: return 8'h76;
         57: return 8'h5b;
         58: return 8'ha2;
         59: return 8'h49;
         60: return 8'h6d;
         61: return 8'h8b;
         62: return 8'hd1;
         63: return 8'h25;
         64: return 8'h72;
         65: return 8'hf8;
         66: return 8'hf6;
         67: return 8'h64;
         68: return 8'h86;
         69: return 8'h68;
         70: return 8'h98;
         71: return 8'h16;
         72: return 8'hd4;
         73: return 8'ha4;
         74: return 8'h5c;
         75: return 8'hcc;
         76: return 8'h5d;
         77: return 8'h65;
         78: return 8'hb6;
         79: return 8'h92;
         80: return 8'h6c;
         81: return 8'h70;
         82: return 8'h48;
         83: return 8'h50;
         84: return 8'hfd;
         85: return 8'hed;
         86: return 8'hb9;
         87: return 8'hda;
         88: return 8'h5e;
         89: return 8'h15;
         90: return 8'h46;
         91: return 8'h57;
         92: return 8'ha7;
         93: return 8'h8d;
         94: return 8'h9d;
         95: return 8'h84;
         96: return 8'h90;
         97: return 8'hd8;
         98: return 8'hab;
         99: return 8'h00;
         100: return 8'h8c;
         101: return 8'hbc;
         102: return 8'hd3;
         103: return 8'h0a;
         104: return 8'hf7;
         105: return 8'he4;
         106: return 8'h58;
         107: return 8'h05;
         108: return 8'hb8;
         109: return 8'hb3;
         110: return 8'h45;
         111: return 8'h06;
         112: return 8'hd0;
         113: return 8'h2c;
         114: return 8'h1e;
         115: return 8'h8f;
         116: return 8'hca;
         117: return 8'h3f;
         118: return 8'h0f;
         119: return 8'h02;
         120: return 8'hc1;
         121: return 8'haf;
         122: return 8'hbd;
         123: return 8'h03;
         124: return 8'h01;
         125: return 8'h13;
         126: return 8'h8a;
         127: return 8'h6b;
         128: return 8'h3a;
         129: return 8'h91;
         130: return 8'h11;
         131: return 8'h41;
         132: return 8'h4f;
         133: return 8'h67;
         134: return 8'hdc;
         135: return 8'hea;
         136: return 8'h97;
         137: return 8'hf2;
         138: return 8'hcf;
         139: return 8'hce;
         140: return 8'hf0;
         141: return 8'hb4;
         142: return 8'he6;
         143: return 8'h73;
         144: return 8'h96;
         145: return 8'hac;
         146: return 8'h74;
         147: return 8'h22;
         148: return 8'he7;
         149: return 8'had;
         150: return 8'h35;
         151: return 8'h85;
         152: return 8'he2;
         153: return 8'hf9;
         154: return 8'h37;
         155: return 8'he8;
         156: return 8'h1c;
         157: return 8'h75;
         158: return 8'hdf;
         159: return 8'h6e;
         160: return 8'h47;
         161: return 8'hf1;
         162: return 8'h1a;
         163: return 8'h71;
         164: return 8'h1d;
         165: return 8'h29;
         166: return 8'hc5;
         167: return 8'h89;
         168: return 8'h6f;
         169: return 8'hb7;
         170: return 8'h62;
         171: return 8'h0e;
         172: return 8'haa;
         173: return 8'h18;
         174: return 8'hbe;
         175: return 8'h1b;
         176: return 8'hfc;
         177: return 8'h56;
         178: return 8'h3e;
         179: return 8'h4b;
         180: return 8'hc6;
         181: return 8'hd2;
         182: return 8'h79;
         183: return 8'h20;
         184: return 8'h9a;
         185: return 8'hdb;
         186: return 8'hc0;
         187: return 8'hfe;
         188: return 8'h78;
         189: return 8'hcd;
         190: return 8'h5a;
         191: return 8'hf4;
         192: return 8'h1f;
         193: return 8'hdd;
         194: return 8'ha8;
         195: return 8'h33;
         196: return 8'h88;
         197: return 8'h07;
         198: return 8'hc7;
         199: return 8'h31;
         200: return 8'hb1;
         201: return 8'h12;
         202: return 8'h10;
         203: return 8'h59;
         204: return 8'h27;
         205: return 8'h80;
         206: return 8'hec;
         207: return 8'h5f;
         208: return 8'h60;
         209: return 8'h51;
         210: return 8'h7f;
         211: return 8'ha9;
         212: return 8'h19;
         213: return 8'hb5;
         214: return 8'h4a;
         215: return 8'h0d;
         216: return 8'h2d;
         217: return 8'he5;
         218: return 8'h7a;
         219: return 8'h9f;
         220: return 8'h93;
         221: return 8'hc9;
         222: return 8'h9c;
         223: return 8'hef;
         224: return 8'ha0;
         225: return 8'he0;
         226: return 8'h3b;
         227: return 8'h4d;
         228: return 8'hae;
         229: return 8'h2a;
         230: return 8'hf5;
         231: return 8'hb0;
         232: return 8'hc8;
         233: return 8'heb;
         234: return 8'hbb;
         235: return 8'h3c;
         236: return 8'h83;
         237: return 8'h53;
         238: return 8'h99;
         239: return 8'h61;
         240: return 8'h17;
         241: return 8'h2b;
         242: return 8'h04;
         243: return 8'h7e;
         244: return 8'hba;
         245: return 8'h77;
         246: return 8'hd6;
         247: return 8'h26;
         248: return 8'he1;
         249: return 8'h69;
         250: return 8'h14;
         251: return 8'h63;
         252: return 8'h55;
         253: return 8'h21;
         254: return 8'h0c;
         255: return 8'h7d;
      endcase;

endmodule
