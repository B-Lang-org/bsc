// Package that defines a synonym using Helper's synonym
// This creates a synonym chain for testing

package HelperAlias;

import Helper::*;

// Synonym that uses Helper's Byte synonym
typedef Byte MyByte;

export MyByte;

endpackage
