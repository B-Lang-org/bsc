function bit[3:0] f();
  bit[3:0] x = 3;
  f = x;
endfunction
