interface Id;
   method a id(a in);
endinterface
