Bool x = True;

Bool y = x[0];

