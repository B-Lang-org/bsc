`define size 2
`define modName sysTest2

`include "Test.bsv"

