String foo;
foo = "foo\n";

