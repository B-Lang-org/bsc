module mkTest1 (Empty);
    Reg#(Int#(32)) x <- mkReg;
endmodule
