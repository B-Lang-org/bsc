// Test that a non clock name is not OK

(* synthesize *)
(* gate_input_clocks="c" *)
module sysGateInputClocks4 #(Clock c1, Clock c2, Clock c3) ();
endmodule
