package ReExportSame_Q;

export T(..);

typedef union tagged {
  Bool Tag1;
  Bool Tag2;
 } T;

endpackage
