Bit #(5) x;
x = 5;
Bit #(7) y;
y = 7;
Bit #(12) z;
z = {x,y};
