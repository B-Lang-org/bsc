package ModuleAugmented() where
{}
