function Bool f();
  for (int x=1, int z=3; x<3; int x, x=x+1)
  begin
    z = z + x;
  end
  return False;
endfunction
