package ReExportPkg_Q (package ReExportPkg_P) where

import ReExportPkg_P

