module mkFoo();
  rule bogus();
  endrule
endmodule
