package IfLifting(sysIfLifting) where

-- Lifting of if-branches: `b.set False' and `b.set True' on two sides
-- of the `if' should be lifted out to `b.set (nosplitIf a False True)'

sysIfLifting :: Module Empty
sysIfLifting =
  module
    a :: Reg Bool
    a <- mkRegU
    b :: Reg Bool
    b <- mkRegU
    rules
        when True ==> (nosplitIf a (b := False) (b := True))

