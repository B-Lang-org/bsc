module mkTest();
  Integer x;
  Bool y;
  { x, y, z } = tuple3(0,True,1);
endmodule

