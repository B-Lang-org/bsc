import Vector::*;

export Vector::*;
export Vector::*;

