(* synthesize *)
(* clock_prefix="foo bar" *)
module sysCLKAttribWithSpace ();
endmodule

