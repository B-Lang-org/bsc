// test generation of undefined values across package boundaries

import HiddenType::*;

(* synthesize *)
module sysPackageTest();
  mkFoo();
endmodule



