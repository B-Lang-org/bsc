package DegreePrimeSymbol((°´), (´°), (+´), (+°)) where

(°´) :: a -> b -> (a, b)
x °´ y = (x,y)

(´°) :: a -> b -> (a, b)
x ´° y = (x,y)

(+´) :: a -> b -> (a, b)
x +´ y = (x,y)

(+°) :: a -> b -> (a, b)
x +° y = (x,y)
