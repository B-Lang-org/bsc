import Vector::*;

(* synthesize *)
module sysRenamePort ( (* port="B" *)Vector#(2,Bool) bs, Empty ifc);
endmodule

