package StructPat_DupField_BothQual where

import FloatingPoint

-- The bad qualifier is on the second field to test that,
-- even though type disambiguation was done using the first field,
-- the qualifiers on later fields are still considered
-- (and reported as an error when they don't match)

fn :: FloatingPoint.Half -> Bool
fn (FloatingPoint.Half { FloatingPoint.sign = True; Foo.sign = b }) = b
fn _ = False
