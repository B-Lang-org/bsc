(* synthesize *)
module mkWrongTop ();
   let m <- mkRightMod;
endmodule

(* synthesize *)
module mkRightMod ();
endmodule

