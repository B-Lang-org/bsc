package ClassWithDefault (C(..)) where

class C a where
  f :: a -> Bool
  g :: a -> Bool
  g x = not (f x)
  h :: a -> Bool
  i :: a -> Bool

-- warn about missing "i" but not "g"
instance C Integer where
  f x = x > 17
  h x = x > 2

v :: Integer
v = 5

-- should use the proper definition of "g"
{-# verilog sysClassWithDefault #-}
sysClassWithDefault :: Module Empty
sysClassWithDefault =
  module
    rules
      "r":
        when True
          ==> action
                if (g v) then $display "1yes" else $display "1no"
                if (f v) then $display "2yes" else $display "2no"

