module sysTwoActions();
   Action a1=action
      int i=16;
      int bad=True;
      $display("Hello ",i);
   endaction;
   Action a2=action
      int j=12;
      int worse=False;
      $display("world ",j);
   endaction;
endmodule
