package ReExportSame_Sub;

import ReExportSame_P::*;

export ReExportSame_P::*;

endpackage

