`include "defs.incl"

