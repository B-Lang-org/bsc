a foo = 1;