
(* synthesize *)
module sysLiteral_Neg();
   Reg#(Bit#(11)) rg <- mkReg(-'h1);
endmodule

