package ClassDefFieldIsNum () where

class Foo a where
    bar :: 12

