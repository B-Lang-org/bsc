`define FOO

`undef

FOO

`ifndef FOO
Bool x = True;
`endif


