package SignatureTooGeneral() where

-- Expect a "Signature too general" error

foo :: a
foo = 1 :: Integer
