import List::*;

List#(Bool) xs = List::nil;
