interface Ifc #(type a, type b, type a);
  method Action m();
endinterface
