(* synthesize *)
(* doc = "This appears twice" *)
(* doc = "This is unique" *)
(* doc = "This appears twice" *)
(* doc = "This is also unique" *)
module sysDuplicateCommentOnModule();
endmodule

