`define size 1
`define modName sysTest1

`include "Test.bsv"

