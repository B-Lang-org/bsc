(* synthesize *)
(* no_default_reset *)
module sysNoDefaultReset_Inout#(Inout#(Bool) io)();
endmodule
