import ConDup_Leaf::*;

// Re-export the same type, but with hidden constructors
export U;

