package Five(five) where

five :: Bool -> Integer
five x = 5

