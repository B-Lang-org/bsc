Integer a = 42;
Integer b = 'd42;
Int#(32) c = 32'd42;
Integer d = 'h2a;
Int#(32) e = 32'h2a;
Integer f = 'o52;
Int#(32) g = 32'o52;
Integer h = 'b101010;
Int#(32) i = 32'b101010;
