
(* synthesize *)
module sysSizedLiteral_Neg();
   Reg#(Bit#(11)) rg <- mkReg(-11'h1);
endmodule

