function Action f(Bool x1, Bool x2, Bool x3);
   $display(x1, x2, x3);
endfunction

Action b = f(False, True, False, True);

