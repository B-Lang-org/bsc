import FieldDup_Leaf::*;

// Re-export the same type, but with hidden fields
export S;

