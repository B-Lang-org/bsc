export Ptak;

typedef union tagged {
   Bool Żuraw;
   void Gżegżółka;
} Ptak;

