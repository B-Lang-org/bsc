// Bug 1336

import "BVI"
   module mkImportModIfc_TooManyArgs(Reg#(Bool,Bool));
      default_clock no_clock;
      default_reset no_reset;
   endmodule

