package Bug437(foo) where

foo :: Integer
foo = True
