typedef union tagged {
} TaggedUnionEmpty;

