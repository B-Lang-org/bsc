Bit#(4) x = 17;
Bit#(3) y = x;

