// Second level include
typedef Bool BBOO ;

`include "IncDep2.bsv"
