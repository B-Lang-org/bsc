int someint;
someint = 1;

Int#(32) otherint;
otherint = someint;
