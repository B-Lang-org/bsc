
Bit#(11) x = 11'h800;

