package TypeAliasResGivenNonNumIsNumParam () where

type (Foo :: # -> *) a = a

