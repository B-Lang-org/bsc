module sysECtxRedIsModuleActionValue_AVExprInModBlock(Empty);
   $display("Hello");
   rule r;
      $display("World");
   endrule
endmodule
