module sysAmbigTCon_TSub (Reg#(Bit#(TSub#(x,y))));
endmodule
