function int f (int n);
  case (n) matches
    0: return 17;
    ._: return (_+1);
  endcase
endfunction
