// Third helper that uses Helper's Color type

package Helper3;

import Helper::*;

function Bool isRed(Helper::Color c);
    return c == Red;
endfunction

export isRed;

endpackage
