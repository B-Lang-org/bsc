
Bit#(11) x = 0'h1;

