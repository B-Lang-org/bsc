Action a1;
a1 = $finish;

Action a2;
a2 = $display;

Action a3;
a3 = $stop;
