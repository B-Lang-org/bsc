package EmptyModule_Layout where

m :: Module Empty
m = module

x :: Integer
x = 17
