module mkBug423_1();
  rule first;
  // endrule (supposedly forgotten)

  rule second;
  endrule
endmodule
