import Vector::*;

(* synthesize *)
module sysRenameReset ( (* reset="R" *)Vector#(2,Reset) rsts, Empty ifc);
endmodule

