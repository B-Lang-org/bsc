package FailIAp where

import BuildVector
import Vector

shuffle :: Vector 4 (Bit 64) -> Vector 4 (Bit 64)
shuffle vs =
    let reordered = fmap ((!!) vs) $ vec 1 2 3 0
    in  reordered
