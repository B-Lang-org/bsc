package VarDefn_NoType () where

_ = True

