package Latin1MultilineComment(foo) where

{-
   comment �
   with � a � non-ASCII
   � symbol
 -}

foo :: (Bits a sza) => a -> a
foo = unpack `compose` pack

