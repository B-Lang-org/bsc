import Prelude::mkReg;
