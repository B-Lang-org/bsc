(*synthesize*)
module connectIntegers#(Inout#(Integer) x, Inout#(Integer) y)();
endmodule
