function Action f();
   $display("foo");
endfunction

Action a = f(True, False, True);

