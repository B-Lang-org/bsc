import "BVI"
module mkBug1470 ();
   port P = 1'b1;
endmodule

