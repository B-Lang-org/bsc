package NonNumWhereNumExpected () where

x :: Bit Bool
x = 0

