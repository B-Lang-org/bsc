module mkFoo();
  id(mkFoo());
endmodule
