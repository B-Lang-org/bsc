package EHasImplicit2(mkPort, mkTop) where

import FIFO

{-# verilog mkPort #-}
mkPort :: Bit 16  -> Module Empty
mkPort x = module 
            rules
             when True ==> action
                            $display x
                            $finish 0

mkTop :: Module Empty
mkTop = module 
          f :: FIFO (Bit 16) <- mkFIFO
          p :: Empty <- mkPort (f.first)

