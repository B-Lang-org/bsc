import "BVI" StringParamErr2 =
module vStringParamErr2#(String s)(Empty ifc);
   port foo = s;

endmodule
