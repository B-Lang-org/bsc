package Zow;


module mkZow (Empty);
   
   Reg#(Bool) zow2 <- mkReg(False);
   
endmodule


endpackage