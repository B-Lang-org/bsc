function int \+ (int a, int b);
  return ?;
endfunction
