import Sub1::*;

(*synthesize*)
module mkTest ((*port="VAL"*)Bool x, Ifc1 i);
endmodule

