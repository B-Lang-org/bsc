
`define m(x

Bool b = `m(True) && True;

Bool b2 = `m(False);
