function bit[3:0] f();
  module mkBogus();
  endmodule
  f = 3;
endfunction

