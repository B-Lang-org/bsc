-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EBitSel.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the EBitSel error of the bluespec
-- compiler (Bit Selection Out of Range)
--
-- Error produced when generating verilog for mkShifter64
-----------------------------------------------------------------------

package EBitSel (Shifter, mkShifter64) where

-- import UInt
import Push
import GetPut
import ClientServer

type Shifter n =
    Server (UInt n {-value-}, UInt (TLog n) {-shift amt-}) (UInt n {-result-})

{-# verilog mkShifter64 #-}
mkShifter64 :: Module (Shifter 64)
mkShifter64 =
    module (getResult, putResult) :: (Get (UInt 64), Put (UInt 64)) <- mkGPFIFO
           shifter :: Push (UInt 64, UInt 6)
                   <- (passed shift1 �
                       passed shift1 �
                       qbuffer �
                       passed shift1 �
                       passed shift1 �
                       qbuffer �
                       passed shift1 �
                       passed shift1 �
                       passed strip �
                       pass � tee (putResult.put) �
                       sink)
           interface
             request = interface Put { put (val,by) = shifter.push (val,by) }
             response = getResult

-- one shift stage
shift1 :: (Add 1 m' m) => (UInt n, UInt m) -> (UInt n, UInt m')
shift1 (val, by) = let i = fromInteger (valueOf m')
                       shift = (pack by)[2:2] == 1
                       val' = if shift then val << (1 << i) else val
                       by' = truncate by
                   in  (val', by')

-- signature ensures that no stages are missing
strip :: (UInt n, UInt 0) -> UInt n
strip (x,_) = x






