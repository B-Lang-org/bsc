package StructDefn_Field () where

struct S =
  _ :: Bool

