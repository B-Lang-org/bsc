export sysStateNameTest2;

(* synthesize *)
module sysStateNameTest2(Empty);
   Reg#(Bit#(16)) b <- mkReg(11);
endmodule 
