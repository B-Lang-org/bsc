
interface Ifc;
 (* ready = "" *)
 method Bool check ();
endinterface

