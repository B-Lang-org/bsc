function Bool f();
  Bool x;
  f = True;
endfunction
