import ReExportItems_P::*;

export AB(..);

export a;
