module sysECtxRedIsModuleActionValue_ModBindInAVBlock();
   rule r;
      let rg <- mkReg(0);
   endrule
endmodule

