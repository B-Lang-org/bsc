interface Bogus#(type a) provisos Arith#(a)
   method a id(a val);
endinterface
