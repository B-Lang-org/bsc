package DeprecatedLibrary where

{-# properties myFunc = { deprecate = "Replaced by myFunc2." } #-}
myFunc :: Bool -> Bool
myFunc = not

