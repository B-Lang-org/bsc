package Joe(sysJoe) where
import List
import FIFO

--import GetPut
class Put c where
    put    :: c a -> a -> Action

class Get c where
    get    :: c a -> a
    drop   :: c a -> Action

instance Put FIFO where
    put f x  = f.enq x

instance Get FIFO where
    get f    = f.first
    drop f   = f.deq

mkJoint :: (Put o, Get i) => o a -> i a -> Module Empty
mkJoint o i =
    module
      rules
	when True
	 ==> action
		put o (get i)
		drop i

join :: (Put o, Get i) => List (i a) -> o a -> Module Empty
join is o =
    module
	mapM (mkJoint o) is
	return $ interface Empty { }

sysJoe :: Module Empty
sysJoe =
    module
	is :: List (FIFO Nat)
	is <- mapM (\ _ -> mkFIFO) (upto 1 3)
	o :: FIFO Nat
	o <- mkFIFO
	join is o
