package LedDecoder (mkLedDecoder, LedDecoder(..), LedDisplay, LedDigit) where

type LedDisplay = Bit 7
type LedDigit = Bit 4

interface LedDecoder =
  decode :: LedDigit -> LedDisplay

mkLedDecoder :: Module LedDecoder
mkLedDecoder =
    return $
	interface LedDecoder
	    decode x = 
	        case x of
		   0x0 -> 0b1110111
		   0x1 -> 0b0010010
		   0x2 -> 0b1011101
		   0x3 -> 0b1011011
		   0x4 -> 0b0111010
		   0x5 -> 0b1101011
		   0x6 -> 0b1101111
		   0x7 -> 0b1010010
		   0x8 -> 0b1111111
		   0x9 -> 0b1111011
		   0xa -> 0b1111110
		   0xb -> 0b0101111
		   0xc -> 0b0001101
		   0xd -> 0b0011111
		   0xe -> 0b1101101
	           0xf -> 0b1101100
