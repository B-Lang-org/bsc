(* synthesize *)
module mkDummyModule(Empty);
endmodule

