function Action f(Bool x1, Integer x2, Bool x3);
   $display(x1, x2, x3);
endfunction

Action a = f(True, False, True);

