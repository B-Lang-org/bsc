package Environment(	) where { }

