function Action f();
  action
    bit[3:0] x = 3;
  endaction
endfunction
