(* synthesize *)
module sysStringHead_Empty();
   rule r;
      $display(stringHead(""));
   endrule
endmodule
