ActionValue#(Bool) av;
av =
  actionvalue
    return id(True);
  endactionvalue;
