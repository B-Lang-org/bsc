package ReExportPkg_Top (x, y, z) where

import ReExportPkg_Q

x :: T
x = 3

-- This should compile (tests "T2" type, "T2" constructor, and value "v")
y :: T2
y = T2 v

-- This should compile
-- (And tests that instances are exported too)
z :: T
z = 2 + x

