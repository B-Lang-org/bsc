function Bool listy();
  Bool xsss[2][3][5][8];
  listy = xsss[0][2][4][6];
endfunction
