package Five(five) where

five :: Bool -> Integer
five x = if x then 5 else 0

