-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EUnify.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the EUnify error of the bluespec
-- compiler
--
-----------------------------------------------------------------------


package EUnify() where

-- import Int

sum :: Int 2 -> Int 2 -> Int 3
sum x y = x + y;



