module mkTest ();
  Tuple3#(Bool, Integer, Bit#(8)) {b,i,v};
  //{b,i,v} = tuple3(True,1,2);
endmodule
