package Latin1Code(foo) where

foo :: (Bits a sza) => a -> a
foo = unpack � pack

