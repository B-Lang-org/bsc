package NoArgPlusOne () where

x :: Bool Bool
x = _

