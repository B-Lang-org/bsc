Bool foo;
foo = True;
Bool bar;
bar = False;
