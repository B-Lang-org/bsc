function Bool listy();
  Bool xsss[2][3][4][5][6][6][5][4][3][2];
  listy = xsss[1][2][3][4][5][5][4][3][2][1];
endfunction
