
interface Ifc;
  (* enable = " name" *)
  method Action start(Bool a, Bool b);
endinterface

