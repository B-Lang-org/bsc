Bool _ = True;

// Test that "_" can be used for Bool
Bool y = ! _;

