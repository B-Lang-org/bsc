(* gate_prefix="", gate_input_clocks="default_clock" *)
module sysEmptyCLKAttrib ();
endmodule

