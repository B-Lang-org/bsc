package OneArgPlusOne () where

x :: Bit 1 2
x = _

