package TLM;

import TLMDefines::*;

export TLMDefines::*;

endpackage
