package Test() where

f :: Bool
f = (1.0 > 0)

