/**** this file tests a multi-line comment

this is junk
**/
package Comment;
Bool x = True;
// Another comment
/* a single-line comment */
/* another multi-line comment

*/
endpackage
