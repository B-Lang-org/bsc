package StructUpd_DupField_QualAndUnqual where

import FloatingPoint

fn :: FloatingPoint.Half -> FloatingPoint.Half
fn x = x { sign = True; FloatingPoint.sign = 0 }
