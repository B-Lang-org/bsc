`define is 500
`define fs 1
`define full sysFromReal_500_1

`include "FromReal.bsv"
