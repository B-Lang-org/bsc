package ReExportPkgBSV_Q;

import ReExportPkg_P::*;

export ReExportPkg_P::*;

endpackage
