module sysExplictActions();
   Action a=True;
   Action b=False;
endmodule
