function Action f();
  action
    bit[3:0] x;
    x = 3;
    x = 7;
  endaction
endfunction
