

import Interfaces :: * ;
import FIFO :: * ;
import FIFOF :: * ;
import GetPut :: * ;
import LFSR :: * ;

interface MasterSlave ;
   interface Master m ;
   interface Slave s ;
endinterface

(* synthesize *)
module mkDMAC( MasterSlave ) ;

   

endmodule
         
