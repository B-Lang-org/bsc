function Bool listy();
  Bool xs[2];
  xs[1] = True;
  listy = xs[0];
endfunction
