typedef union tagged {
  function a id(a in) MyId;
} Id;

