
function Bit#(n) fn();
  return pack(0);
endfunction

