package Defl_NoType () where

x :: Bool
x = let _ = True
    in  True

