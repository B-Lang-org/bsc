
function Reg#(Bool) mkFn();
  return (
     interface Reg;
        Bool x = True;
     endinterface
   );
endfunction

