// Comment

`line(/file/path