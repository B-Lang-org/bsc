-----------------------------------------------------------------------
-- Project: Bluespec

-- File: ENotField1.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers an (ENotField) error

-- Error Message : bsc ENotField1.bs
-- bsc: Compilation errors:
-- "ENotField1.bs", line 51, column 12, Field "result" is not in "ENotField1.ENotField1"
-----------------------------------------------------------------------

package ENotField1 (ENotField1(..), mkENotField1) where

-- import Int

interface ENotField1 =
    start   :: Int 32 -> Int 32 -> Action
    product :: Int 32


mkENotField1 :: Module ENotField1
mkENotField1 =
    module

        x :: Reg (Int 32)
        x <- mkReg 0

	y :: Reg (Int 32)
	y <- mkReg 0

        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0
