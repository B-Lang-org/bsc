
`undef -

Bool x = True;

