package Lambda_Arg () where

x :: Bool
x = (\ _ -> True) False

