package LFSRExtra where

import LFSR
import Vector

import Rules
import VectorExtra

mkAutoStepLFSR :: (IsModule m c, Bits t t_sz) => m (LFSR (Bit t_sz)) -> m t
mkAutoStepLFSR mk = module
  _lfsr :: LFSR (Bit t_sz) <- mk
  always "AutoStepLFSR" _lfsr.next
  return $ unpack _lfsr.value

-- Class to store polynomial values for LFSRs. The polynomials below were taken
-- from three sources. The lfsrPolyK (K for Koopman) values are from first entry
-- of each file in:
--   http://users.ece.cmu.edu/~koopman/lfsr/
-- The lfsrPolyX (X for Xilinx) values are from the Xilinx documentation at:
--   https://docs.xilinx.com/v/u/en-US/xapp052
-- The lfsrPolyC (C for Computed) values are computed using modified code from:
--   http://www.seanerikoconnor.freeservers.com/Mathematics/AbstractAlgebra/PrimitivePolynomials/overview.html
-- Note: The K ones are probably best to use where possible, since they are the
-- ones used in LFSR.bs, and they tend to include taps at the low end of the
-- register, which will produce sequences which initially contain more nonzero
-- bits on the low end. But, there are 168 of the X ones, and only 64 of the K
-- ones. Regardless, the issue with starting with many 0s can be avoided by
-- using a seed. The C ones appear to be similar to the K ones, but they can be
-- computed and added to this file as we need more.

class LFSR_Polys n where
  lfsrPolyK :: Maybe (Bit n)  -- K for Koopman
  lfsrPolyK = Invalid
  lfsrPolyX :: Maybe (Bit n)  -- X for Xilinx
  lfsrPolyX = Invalid
  lfsrPolyC :: Maybe (Bit n)  -- C for Computed
  lfsrPolyC = Invalid

-- Select a polynomial to use for the LFSR. Prefer K where possible.
lfsrPoly  :: (LFSR_Polys n) => Bit n
lfsrPoly = case (lfsrPolyK, lfsrPolyX, lfsrPolyC) of
  (Valid k, _, _)             -> k  -- Prefer K where possible.
  (Invalid, Valid x, _)       -> x  -- Fall back to X.
  (Invalid, Invalid, Valid c) -> c  -- Fall back to C.
  (Invalid, Invalid, Invalid) -> error "No LFSR polynomial for this size."

-- Similar to mkFeedLFSR, but with a seed value.
mkLFSRSeed :: (IsModule m c, LFSR_Polys n) => Bit n -> m (LFSR (Bit n))
mkLFSRSeed s = module
  r :: Reg (Bit n) <- mkRegA s
  interface
    seed  = r._write
    value = r
    next  = r := let lsb = r[0:0]
                     sh = r >> 1
                     x  = if lsb == 1 then lfsrPoly else 0
                  in sh ^ x

-- Use seed = 1 by default, since that is what mkFeedLFSR uses in LFSR.bs.
mkLFSR :: (IsModule m c, LFSR_Polys n) => m (LFSR (Bit n))
mkLFSR = mkLFSRSeed 1

type LFSRSeedLen = 928  -- The longest LFSR that is currently available.
type NumLFSRSeeds = 17  -- The number of seeds that are available.

-- Note: It is important that each seed be nonzero regardless of how it is
-- truncated. If an LFSR is created with an all-zero seed, it will only ever
-- produce 0s. So, the low bit is explicitly set, and the rest are "random".
-- from python:   hex(secrets.randbits(...) | 1)
-- http://xkcd.com/221

lfsrSeeds :: Vector NumLFSRSeeds (Bit LFSRSeedLen)
lfsrSeeds = vec
  0x1bca484aeebc0e9c7bb9dda5e4dd7c3061635ae2bd45b09d0d98fd0d1d9c6db9aa85ac764c6a15928316d2e0ecc2c61195212d27d7ffa70ff17cba62e9a346d74a9db6377897218eb69ca8b95298f9022220a4c528a7abb4b43417e3e56dd3557cdef08d702e66eb5837a8cb8f6a4e21efb663c5
  0xd3d4a023c7c49ccffb8301242f33c9ef62873f113cc540fc81e53b03e9c84993705fe134ffa6f0a0c8ee3d77eca6a7f8059dba7b759c5c4ca374fc308d4183ebdbe836bc3f9b5c40dc0ea9b852aa250357aa51746b060d3d32a359739cfb1c1882a2994cc6f6a67b41e3f69d5e12c5fcdb0eb4b9
  0x3ddebb0a6013de1aae1d7662fa502e8440def108a3456efa35e03e6a078595e2a65089971aad07741c59ea17eb0bb198bdd8e4778c6fa8c5930536ee4202fd20ae2bf68134f8d60da080685898f6e917ca0cb8b539c2907480fec94145c50bdf6170bb96eb5e9048e5145d1d8a8209ab31735049
  0xc935f9706ed50cb2dc50e13a9520ef747c8c9655db062bb6bf78de72820f6bf2f19394fb40adff2beeec39be8e861848f7b39b0123b8f585bf38d552d7e96716ff3c84ffd65e736c563a18a0e01c707cf6f9ab0e8aebbff0cfc2d3df5320f6a6ecba0367015884cb82b00e915ea072365456415f
  0xee1d9f70a02584172aedeaf5f7a4e0a6a65cee3935ad2ad550ebc74975a45c19a366973d0e148b893001a1150a1c13ba42f43c472d1a788c79487e78ab684b05a0aef477b6057ce794a9d5529fc94f15208d27b8cd754170ed84e3a38ebf7199708cec4226f3d32fc528a65006323ecd250e70e9
  0xa17d29113e5d0e4ebb223d1285a74dccd8d2f340397081bd4de6e6dafee4150a577b8d6db4954ba4452a5651446e44dfb421f875649fbb6719fdc5428c850845491807ccb9e7bbcf94bcf848e9bd1699b7a647bab2fd11f57f5f64b08f04795aab4560427bc30e8379211bb7d112ae23c50da509
  0x84ae2c72fee933acb98f6dff0a3d691745c2f5579648d1abfc20528aa4b6ff2f7a660945ac635af05ef04596062b38ae9521977e518391b1fd10ccd902c0d300c555ae125231a403b4ab27e6d482e951a0d03e232f07dd3547e03e80d6535d0debfea882cb423768f427ee4cc7941439fa2a0f39
  0x4644725977ab4c704ae8325c8ef4335d399e0b594bf78d8a79f893cb9fcf481cba3a0b4b388b3d4fe871d6a791f9fa120190cb4887d8b3e5ffe693b6043ee0e1c06ae53cdd6f47befb1dfd4a0fe02aa845d5057d4afddb09fdfd8d9168fbf95af022da4c729600a7b750196d523ace581d006ec9
  0x2aa345f73206d3bdf15a2ed720af978c8ab48211b204a1e8b23c79463608fabb5fc9d99d053f10dd86e8f96d2fd7daadbbf945d3e5e75992196fd4f849c53109a7f400969be39ae7c7e811488406a2c55febeece84f48754c29e0c188783a42875e12277e7ed7710d0d4845178ac09178e3ba71b
  0x53440a0eb5d43040b854d416c571c2b770b3e8575af6cbd27ab6b326522401b6ee54a5499cab461cc92f7b9ff5bada9b6cee014ce9d13f4cb1d72a23b7175518a737e3211db9b2140fe72f8ff72bd02c96553f07cf8f40f167730035cd426515296b415c6f022c08edcf6f434b8e1513dac65b21
  0x3dc6b9e6e866b918ed8277382870c13f7f5a1c92c2ca88340f8a0b9750608a96e40676ed79037aef99cc08f720e6110fb2ca68f382eeebc254d22b06d90eb076536e545689e8e2408f2b90aadd34334a397e1dd079f06f54c92f5089d63c2086e29f663d7d5501dd023c4510adb73eeccf0fd95d
  0xeb422e445fcec69a10ac630f71e73e3cf2fde2efce85f1c967933d9aa9358cede98bf288922e72e52934fdd02a0fdc57398e26ebab501eebe058026790128cb6bc0f22a9306e7a1eeeec142f18193a30adc68336875fe5e3754095ba122b755187a976b4e952decb03a049bb9f2706dd836e2f8f
  0x44ea77d14880e90f8a84ad67398567aa6c6be48596d715e0e6c0880caef59cfb14a0212703ab251ecf3be83dc06b7185c8614556004364275f860c82b993ac9032565fe7565697ebf4f5879e61b48144b685c9caf048995526c3f13bbe5c593fb0152f8858321e61f5b636a5ce076377749da45f
  0x26ab168536cbe68bd71c07ed79d014d56619a2fe8f11144e6d8cf262428f9290b97845d2e024c133d3c08da10215b43601514d85365fe342b5cf56b355fe0b3cb618ff2842d19867df6199375e82f9530f88cf8718e948c3c461304f3028172fa6c40f4fe7c44f94723c8dc3dc396710c0b746dd
  0xcb81008e510b2a992c3056b2b383f0065f971240f5728732a3f3642af5bfdaa78bbcf0178998b9c94411420433b000bc78075571fbb6a21920d1ea2ec468a8405e1345aedea95d57fdee1c667397df3ea20ced718c223d082a16709cd15453f97d063a853070902f83cd44b8668e71b984b97127
  0xacfd199c88e44b06a1a9c7933e2c687034f5aafbebf26275718ab02035216847fb1054ffdf65ebb249de6c605877b47baa43add24a9639cc3d3451e5184002c15078f1323924119b3711bd932bbe80b86f308e794e02ac2db75575191320b6e5c09f8bc202d594a66ca9dba45735d3a0fb786d37
  0xcb2869d20885ad4a191a6259dba61af3e4a04103abcffe7b81c68c83ef14a6ef3b88d9431779a130b4ede6225fb2455468652a514083619eff5cfc6dc1a29faff60ca19a2c37699837c972ebc69b102b3f4c1715c153e11e5954487204512707a95a6fe065bed7a02ff80971424982eea4b15c8d

-- For cases where a seed that isn't "mostly 0s" is desired. The integer is just
-- a seed to make it easy to generate some seeded LFSRs that start with
-- different values.
mkLFSRRandSeedN :: (IsModule m c, LFSR_Polys n, Add p n LFSRSeedLen) =>
  Integer -> m (LFSR (Bit n))
mkLFSRRandSeedN i = mkLFSRSeed $ truncate $
  lfsrSeeds !! (((valueOf n) + i) % (valueOf NumLFSRSeeds))

mkLFSRRandSeed :: (IsModule m c, LFSR_Polys n, Add p n LFSRSeedLen) =>
  m (LFSR (Bit n))
mkLFSRRandSeed = mkLFSRRandSeedN 0

-- All the LFSR polynomials:
instance LFSR_Polys 2 where
  lfsrPolyX = Valid 0x3  -- This one was actually taken from the Wikipedia page.
  lfsrPolyC = Valid 0x3
instance LFSR_Polys 3 where
  lfsrPolyX = Valid 0x6
  lfsrPolyC = Valid 0x5
instance LFSR_Polys 4 where
  lfsrPolyK = Valid 0x9
  lfsrPolyX = Valid 0xc
  lfsrPolyC = Valid 0x9
instance LFSR_Polys 5 where
  lfsrPolyK = Valid 0x12
  lfsrPolyX = Valid 0x14
  lfsrPolyC = Valid 0x12
instance LFSR_Polys 6 where
  lfsrPolyK = Valid 0x21
  lfsrPolyX = Valid 0x30
  lfsrPolyC = Valid 0x21
instance LFSR_Polys 7 where
  lfsrPolyK = Valid 0x41
  lfsrPolyX = Valid 0x60
  lfsrPolyC = Valid 0x41
instance LFSR_Polys 8 where
  lfsrPolyK = Valid 0x8E
  lfsrPolyX = Valid 0xb8
  lfsrPolyC = Valid 0x8e
instance LFSR_Polys 9 where
  lfsrPolyK = Valid 0x108
  lfsrPolyX = Valid 0x110
  lfsrPolyC = Valid 0x108
instance LFSR_Polys 10 where
  lfsrPolyK = Valid 0x204
  lfsrPolyX = Valid 0x240
  lfsrPolyC = Valid 0x204
instance LFSR_Polys 11 where
  lfsrPolyK = Valid 0x402
  lfsrPolyX = Valid 0x500
  lfsrPolyC = Valid 0x402
instance LFSR_Polys 12 where
  lfsrPolyK = Valid 0x829
  lfsrPolyX = Valid 0x829
  lfsrPolyC = Valid 0x829
instance LFSR_Polys 13 where
  lfsrPolyK = Valid 0x100D
  lfsrPolyX = Valid 0x100d
  lfsrPolyC = Valid 0x100d
instance LFSR_Polys 14 where
  lfsrPolyK = Valid 0x2015
  lfsrPolyX = Valid 0x2015
  lfsrPolyC = Valid 0x2015
instance LFSR_Polys 15 where
  lfsrPolyK = Valid 0x4001
  lfsrPolyX = Valid 0x6000
  lfsrPolyC = Valid 0x4001
instance LFSR_Polys 16 where
  lfsrPolyK = Valid 0x8016
  lfsrPolyX = Valid 0xd008
  lfsrPolyC = Valid 0x8016
instance LFSR_Polys 17 where
  lfsrPolyK = Valid 0x10004
  lfsrPolyX = Valid 0x12000
  lfsrPolyC = Valid 0x10004
instance LFSR_Polys 18 where
  lfsrPolyK = Valid 0x20013
  lfsrPolyX = Valid 0x20400
  lfsrPolyC = Valid 0x20013
instance LFSR_Polys 19 where
  lfsrPolyK = Valid 0x40013
  lfsrPolyX = Valid 0x40023
  lfsrPolyC = Valid 0x40013
instance LFSR_Polys 20 where
  lfsrPolyK = Valid 0x80004
  lfsrPolyX = Valid 0x90000
  lfsrPolyC = Valid 0x80004
instance LFSR_Polys 21 where
  lfsrPolyK = Valid 0x100002
  lfsrPolyX = Valid 0x140000
  lfsrPolyC = Valid 0x100002
instance LFSR_Polys 22 where
  lfsrPolyK = Valid 0x200001
  lfsrPolyX = Valid 0x300000
  lfsrPolyC = Valid 0x200001
instance LFSR_Polys 23 where
  lfsrPolyK = Valid 0x400010
  lfsrPolyX = Valid 0x420000
  lfsrPolyC = Valid 0x400010
instance LFSR_Polys 24 where
  lfsrPolyK = Valid 0x80000D
  lfsrPolyX = Valid 0xe10000
  lfsrPolyC = Valid 0x80000d
instance LFSR_Polys 25 where
  lfsrPolyK = Valid 0x1000004
  lfsrPolyX = Valid 0x1200000
  lfsrPolyC = Valid 0x1000004
instance LFSR_Polys 26 where
  lfsrPolyK = Valid 0x2000023
  lfsrPolyX = Valid 0x2000023
  lfsrPolyC = Valid 0x2000023
instance LFSR_Polys 27 where
  lfsrPolyK = Valid 0x4000013
  lfsrPolyX = Valid 0x4000013
  lfsrPolyC = Valid 0x4000013
instance LFSR_Polys 28 where
  lfsrPolyK = Valid 0x8000004
  lfsrPolyX = Valid 0x9000000
  lfsrPolyC = Valid 0x8000004
instance LFSR_Polys 29 where
  lfsrPolyK = Valid 0x10000002
  lfsrPolyX = Valid 0x14000000
  lfsrPolyC = Valid 0x10000002
instance LFSR_Polys 30 where
  lfsrPolyK = Valid 0x20000029
  lfsrPolyX = Valid 0x20000029
  lfsrPolyC = Valid 0x20000029
instance LFSR_Polys 31 where
  lfsrPolyK = Valid 0x40000004
  lfsrPolyX = Valid 0x48000000
  lfsrPolyC = Valid 0x40000004
instance LFSR_Polys 32 where
  lfsrPolyK = Valid 0x80000057
  lfsrPolyX = Valid 0x80200003
  lfsrPolyC = Valid 0x80000057
instance LFSR_Polys 33 where
  lfsrPolyK = Valid 0x100000029
  lfsrPolyX = Valid 0x100080000
  lfsrPolyC = Valid 0x100000029
instance LFSR_Polys 34 where
  lfsrPolyK = Valid 0x200000073
  lfsrPolyX = Valid 0x204000003
  lfsrPolyC = Valid 0x200000073
instance LFSR_Polys 35 where
  lfsrPolyK = Valid 0x400000002
  lfsrPolyX = Valid 0x500000000
  lfsrPolyC = Valid 0x400000002
instance LFSR_Polys 36 where
  lfsrPolyK = Valid 0x80000003B
  lfsrPolyX = Valid 0x801000000
  lfsrPolyC = Valid 0x80000003b
instance LFSR_Polys 37 where
  lfsrPolyK = Valid 0x100000001F
  lfsrPolyX = Valid 0x100000001f
  lfsrPolyC = Valid 0x100000001f
instance LFSR_Polys 38 where
  lfsrPolyK = Valid 0x2000000031
  lfsrPolyX = Valid 0x2000000031
  lfsrPolyC = Valid 0x2000000031
instance LFSR_Polys 39 where
  lfsrPolyK = Valid 0x4000000008
  lfsrPolyX = Valid 0x4400000000
  lfsrPolyC = Valid 0x4000000008
instance LFSR_Polys 40 where
  lfsrPolyK = Valid 0x800000001C
  lfsrPolyX = Valid 0xa000140000
  lfsrPolyC = Valid 0x800000001c
instance LFSR_Polys 41 where
  lfsrPolyK = Valid 0x10000000004
  lfsrPolyX = Valid 0x12000000000
  lfsrPolyC = Valid 0x10000000004
instance LFSR_Polys 42 where
  lfsrPolyK = Valid 0x2000000001F
  lfsrPolyX = Valid 0x300000c0000
  lfsrPolyC = Valid 0x2000000001f
instance LFSR_Polys 43 where
  lfsrPolyK = Valid 0x4000000002C
  lfsrPolyX = Valid 0x63000000000
  lfsrPolyC = Valid 0x4000000002c
instance LFSR_Polys 44 where
  lfsrPolyK = Valid 0x80000000032
  lfsrPolyX = Valid 0xc0000030000
  lfsrPolyC = Valid 0x80000000032
instance LFSR_Polys 45 where
  lfsrPolyK = Valid 0x10000000000D
  lfsrPolyX = Valid 0x1b0000000000
  lfsrPolyC = Valid 0x10000000000d
instance LFSR_Polys 46 where
  lfsrPolyK = Valid 0x200000000097
  lfsrPolyX = Valid 0x300003000000
  lfsrPolyC = Valid 0x200000000097
instance LFSR_Polys 47 where
  lfsrPolyK = Valid 0x400000000010
  lfsrPolyX = Valid 0x420000000000
  lfsrPolyC = Valid 0x400000000010
instance LFSR_Polys 48 where
  lfsrPolyK = Valid 0x80000000005B
  lfsrPolyX = Valid 0xc00000180000
  lfsrPolyC = Valid 0x80000000005b
instance LFSR_Polys 49 where
  lfsrPolyK = Valid 0x1000000000038
  lfsrPolyX = Valid 0x1008000000000
  lfsrPolyC = Valid 0x1000000000038
instance LFSR_Polys 50 where
  lfsrPolyK = Valid 0x200000000000E
  lfsrPolyX = Valid 0x3000000c00000
  lfsrPolyC = Valid 0x200000000000e
instance LFSR_Polys 51 where
  lfsrPolyK = Valid 0x4000000000025
  lfsrPolyX = Valid 0x6000c00000000
  lfsrPolyC = Valid 0x4000000000025
instance LFSR_Polys 52 where
  lfsrPolyK = Valid 0x8000000000004
  lfsrPolyX = Valid 0x9000000000000
  lfsrPolyC = Valid 0x8000000000004
instance LFSR_Polys 53 where
  lfsrPolyK = Valid 0x10000000000023
  lfsrPolyX = Valid 0x18003000000000
  lfsrPolyC = Valid 0x10000000000023
instance LFSR_Polys 54 where
  lfsrPolyK = Valid 0x2000000000003E
  lfsrPolyX = Valid 0x30000000030000
  lfsrPolyC = Valid 0x2000000000003e
instance LFSR_Polys 55 where
  lfsrPolyK = Valid 0x40000000000023
  lfsrPolyX = Valid 0x40000040000000
  lfsrPolyC = Valid 0x40000000000023
instance LFSR_Polys 56 where
  lfsrPolyK = Valid 0x8000000000004A
  lfsrPolyX = Valid 0xc0000600000000
  lfsrPolyC = Valid 0x8000000000004a
instance LFSR_Polys 57 where
  lfsrPolyK = Valid 0x100000000000016
  lfsrPolyX = Valid 0x102000000000000
  lfsrPolyC = Valid 0x100000000000016
instance LFSR_Polys 58 where
  lfsrPolyK = Valid 0x200000000000031
  lfsrPolyX = Valid 0x200004000000000
  lfsrPolyC = Valid 0x200000000000031
instance LFSR_Polys 59 where
  lfsrPolyK = Valid 0x40000000000003D
  lfsrPolyX = Valid 0x600003000000000
  lfsrPolyC = Valid 0x40000000000003d
instance LFSR_Polys 60 where
  lfsrPolyK = Valid 0x800000000000001
  lfsrPolyX = Valid 0xc00000000000000
  lfsrPolyC = Valid 0x800000000000001
instance LFSR_Polys 61 where
  lfsrPolyK = Valid 0x1000000000000013
  lfsrPolyX = Valid 0x1800300000000000
  lfsrPolyC = Valid 0x1000000000000013
instance LFSR_Polys 62 where
  lfsrPolyK = Valid 0x2000000000000034
  lfsrPolyX = Valid 0x3000000000000030
  lfsrPolyC = Valid 0x2000000000000034
instance LFSR_Polys 63 where
  lfsrPolyK = Valid 0x4000000000000001
  lfsrPolyX = Valid 0x6000000000000000
  lfsrPolyC = Valid 0x4000000000000001
instance LFSR_Polys 64 where
  lfsrPolyK = Valid 0x800000000000000D
  lfsrPolyX = Valid 0xd800000000000000
  lfsrPolyC = Valid 0x800000000000000d
instance LFSR_Polys 65 where
  lfsrPolyX = Valid 0x10000400000000000
  lfsrPolyC = Valid 0x1000000000000000d
instance LFSR_Polys 66 where
  lfsrPolyX = Valid 0x30180000000000000
  lfsrPolyC = Valid 0x200000000000000b6
instance LFSR_Polys 67 where
  lfsrPolyX = Valid 0x60300000000000000
  lfsrPolyC = Valid 0x40000000000000013
instance LFSR_Polys 68 where
  lfsrPolyX = Valid 0x80400000000000000
  lfsrPolyC = Valid 0x80000000000000051
instance LFSR_Polys 69 where
  lfsrPolyX = Valid 0x140000028000000000
  lfsrPolyC = Valid 0x100000000000000032
instance LFSR_Polys 70 where
  lfsrPolyX = Valid 0x300060000000000000
  lfsrPolyC = Valid 0x200000000000000015
instance LFSR_Polys 71 where
  lfsrPolyX = Valid 0x410000000000000000
  lfsrPolyC = Valid 0x400000000000000015
instance LFSR_Polys 72 where
  lfsrPolyX = Valid 0x820000000001040000
  lfsrPolyC = Valid 0x80000000000000002f
instance LFSR_Polys 73 where
  lfsrPolyX = Valid 0x1000000800000000000
  lfsrPolyC = Valid 0x100000000000000000e
instance LFSR_Polys 74 where
  lfsrPolyX = Valid 0x3000600000000000000
  lfsrPolyC = Valid 0x200000000000000004c
instance LFSR_Polys 75 where
  lfsrPolyX = Valid 0x6018000000000000000
  lfsrPolyC = Valid 0x4000000000000000025
instance LFSR_Polys 76 where
  lfsrPolyX = Valid 0xc000000018000000000
  lfsrPolyC = Valid 0x800000000000000001a
instance LFSR_Polys 77 where
  lfsrPolyX = Valid 0x18000000600000000000
  lfsrPolyC = Valid 0x10000000000000000032
instance LFSR_Polys 78 where
  lfsrPolyX = Valid 0x30000600000000000000
  lfsrPolyC = Valid 0x20000000000000000043
instance LFSR_Polys 79 where
  lfsrPolyX = Valid 0x40200000000000000000
  lfsrPolyC = Valid 0x4000000000000000000e
instance LFSR_Polys 80 where
  lfsrPolyX = Valid 0xc0000000060000000000
  lfsrPolyC = Valid 0x80000000000000000057
instance LFSR_Polys 81 where
  lfsrPolyX = Valid 0x110000000000000000000
  lfsrPolyC = Valid 0x100000000000000000008
instance LFSR_Polys 82 where
  lfsrPolyX = Valid 0x240000000480000000000
  lfsrPolyC = Valid 0x2000000000000000000e9
instance LFSR_Polys 83 where
  lfsrPolyX = Valid 0x600000000003000000000
  lfsrPolyC = Valid 0x40000000000000000004a
instance LFSR_Polys 84 where
  lfsrPolyX = Valid 0x800400000000000000000
  lfsrPolyC = Valid 0x8000000000000000000d5
instance LFSR_Polys 85 where
  lfsrPolyX = Valid 0x1800000300000000000000
  lfsrPolyC = Valid 0x1000000000000000000083
instance LFSR_Polys 86 where
  lfsrPolyX = Valid 0x3003000000000000000000
  lfsrPolyC = Valid 0x2000000000000000000032
instance LFSR_Polys 87 where
  lfsrPolyX = Valid 0x4002000000000000000000
  lfsrPolyC = Valid 0x4000000000000000000051
instance LFSR_Polys 88 where
  lfsrPolyX = Valid 0xc000000000000000018000
  lfsrPolyC = Valid 0x800000000000000000009d
instance LFSR_Polys 89 where
  lfsrPolyX = Valid 0x10000000004000000000000
  lfsrPolyC = Valid 0x10000000000000000000034
instance LFSR_Polys 90 where
  lfsrPolyX = Valid 0x30000c00000000000000000
  lfsrPolyC = Valid 0x20000000000000000000016
instance LFSR_Polys 91 where
  lfsrPolyX = Valid 0x600000000000000000000c0
  lfsrPolyC = Valid 0x40000000000000000000076
instance LFSR_Polys 92 where
  lfsrPolyX = Valid 0xc00c0000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000032
instance LFSR_Polys 93 where
  lfsrPolyX = Valid 0x140000000000000000000000
  lfsrPolyC = Valid 0x100000000000000000000002
instance LFSR_Polys 94 where
  lfsrPolyX = Valid 0x200001000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000031
instance LFSR_Polys 95 where
  lfsrPolyX = Valid 0x400800000000000000000000
  lfsrPolyC = Valid 0x40000000000000000000003b
instance LFSR_Polys 96 where
  lfsrPolyX = Valid 0xa00000000001400000000000
  lfsrPolyC = Valid 0x80000000000000000000006e
instance LFSR_Polys 97 where
  lfsrPolyX = Valid 0x1040000000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000020
instance LFSR_Polys 98 where
  lfsrPolyX = Valid 0x2004000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000004f
instance LFSR_Polys 99 where
  lfsrPolyX = Valid 0x5000000000028000000000000
  lfsrPolyC = Valid 0x4000000000000000000000058
instance LFSR_Polys 100 where
  lfsrPolyX = Valid 0x8000000004000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000c2
instance LFSR_Polys 101 where
  lfsrPolyX = Valid 0x18600000000000000000000000
  lfsrPolyC = Valid 0x10000000000000000000000061
instance LFSR_Polys 102 where
  lfsrPolyX = Valid 0x30000000000000000c00000000
  lfsrPolyC = Valid 0x20000000000000000000000034
instance LFSR_Polys 103 where
  lfsrPolyX = Valid 0x40200000000000000000000000
  lfsrPolyC = Valid 0x4000000000000000000000005e
instance LFSR_Polys 104 where
  lfsrPolyX = Valid 0xc0300000000000000000000000
  lfsrPolyC = Valid 0x800000000000000000000001be
instance LFSR_Polys 105 where
  lfsrPolyX = Valid 0x100010000000000000000000000
  lfsrPolyC = Valid 0x10000000000000000000000003b
instance LFSR_Polys 106 where
  lfsrPolyX = Valid 0x200040000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000031
instance LFSR_Polys 107 where
  lfsrPolyX = Valid 0x5000000000000000a0000000000
  lfsrPolyC = Valid 0x400000000000000000000000057
instance LFSR_Polys 108 where
  lfsrPolyX = Valid 0x800000010000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000037f
instance LFSR_Polys 109 where
  lfsrPolyX = Valid 0x1860000000000000000000000000
  lfsrPolyC = Valid 0x100000000000000000000000001a
instance LFSR_Polys 110 where
  lfsrPolyX = Valid 0x3003000000000000000000000000
  lfsrPolyC = Valid 0x2000000000000000000000000029
instance LFSR_Polys 111 where
  lfsrPolyX = Valid 0x4010000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000004a
instance LFSR_Polys 112 where
  lfsrPolyX = Valid 0xa000000000140000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000000a7
instance LFSR_Polys 113 where
  lfsrPolyX = Valid 0x10080000000000000000000000000
  lfsrPolyC = Valid 0x10000000000000000000000000016
instance LFSR_Polys 114 where
  lfsrPolyX = Valid 0x30000000000000000000180000000
  lfsrPolyC = Valid 0x200000000000000000000000000e6
instance LFSR_Polys 115 where
  lfsrPolyX = Valid 0x60018000000000000000000000000
  lfsrPolyC = Valid 0x40000000000000000000000000057
instance LFSR_Polys 116 where
  lfsrPolyX = Valid 0xc0000000000000000300000000000
  lfsrPolyC = Valid 0x80000000000000000000000000032
instance LFSR_Polys 117 where
  lfsrPolyX = Valid 0x140005000000000000000000000000
  lfsrPolyC = Valid 0x100000000000000000000000000013
instance LFSR_Polys 118 where
  lfsrPolyX = Valid 0x200000001000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000032
instance LFSR_Polys 119 where
  lfsrPolyX = Valid 0x404000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000080
instance LFSR_Polys 120 where
  lfsrPolyX = Valid 0x810000000000000000000000000102
  lfsrPolyC = Valid 0x800000000000000000000000000073
instance LFSR_Polys 121 where
  lfsrPolyX = Valid 0x1000040000000000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000091
instance LFSR_Polys 122 where
  lfsrPolyX = Valid 0x3000000000000006000000000000000
  lfsrPolyC = Valid 0x2000000000000000000000000000023
instance LFSR_Polys 123 where
  lfsrPolyX = Valid 0x5000000000000000000000000000000
  lfsrPolyC = Valid 0x4000000000000000000000000000002
instance LFSR_Polys 124 where
  lfsrPolyX = Valid 0x8000000004000000000000000000000
  lfsrPolyC = Valid 0x8000000000000000000000000000070
instance LFSR_Polys 125 where
  lfsrPolyX = Valid 0x18000000000000000000000000030000
  lfsrPolyC = Valid 0x10000000000000000000000000000057
instance LFSR_Polys 126 where
  lfsrPolyX = Valid 0x30000000030000000000000000000000
  lfsrPolyC = Valid 0x2000000000000000000000000000004a
instance LFSR_Polys 127 where
  lfsrPolyX = Valid 0x60000000000000000000000000000000
  lfsrPolyC = Valid 0x40000000000000000000000000000001
instance LFSR_Polys 128 where
  lfsrPolyX = Valid 0xa0000014000000000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000000000043
instance LFSR_Polys 129 where
  lfsrPolyX = Valid 0x108000000000000000000000000000000
  lfsrPolyC = Valid 0x100000000000000000000000000000010
instance LFSR_Polys 130 where
  lfsrPolyX = Valid 0x240000000000000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000000004
instance LFSR_Polys 131 where
  lfsrPolyX = Valid 0x600000000000c00000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000079
instance LFSR_Polys 132 where
  lfsrPolyX = Valid 0x800000040000000000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000000000003e
instance LFSR_Polys 133 where
  lfsrPolyX = Valid 0x1800000000000300000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000000037
instance LFSR_Polys 134 where
  lfsrPolyX = Valid 0x2000000000000010000000000000000000
  lfsrPolyC = Valid 0x2000000000000000000000000000000051
instance LFSR_Polys 135 where
  lfsrPolyX = Valid 0x4008000000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000002c
instance LFSR_Polys 136 where
  lfsrPolyX = Valid 0xc000000000000000000000000000000600
  lfsrPolyC = Valid 0x8000000000000000000000000000000086
instance LFSR_Polys 137 where
  lfsrPolyX = Valid 0x10000080000000000000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000000009e
instance LFSR_Polys 138 where
  lfsrPolyX = Valid 0x30600000000000000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000000000b6
instance LFSR_Polys 139 where
  lfsrPolyX = Valid 0x4a400000000000000000000000000000000
  lfsrPolyC = Valid 0x40000000000000000000000000000000057
instance LFSR_Polys 140 where
  lfsrPolyX = Valid 0x80000004000000000000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000000000000089
instance LFSR_Polys 141 where
  lfsrPolyX = Valid 0x180000003000000000000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000000000d5
instance LFSR_Polys 142 where
  lfsrPolyX = Valid 0x200001000000000000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000000000079
instance LFSR_Polys 143 where
  lfsrPolyX = Valid 0x600006000000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000000016
instance LFSR_Polys 144 where
  lfsrPolyX = Valid 0xc00000000000000006000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000000000000004a
instance LFSR_Polys 145 where
  lfsrPolyX = Valid 0x1000000000000100000000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000000000031
instance LFSR_Polys 146 where
  lfsrPolyX = Valid 0x3000000000000006000000000000000000000
  lfsrPolyC = Valid 0x2000000000000000000000000000000000016
instance LFSR_Polys 147 where
  lfsrPolyX = Valid 0x6000000003000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000000001f
instance LFSR_Polys 148 where
  lfsrPolyX = Valid 0x8000001000000000000000000000000000000
  lfsrPolyC = Valid 0x8000000000000000000000000000000000054
instance LFSR_Polys 149 where
  lfsrPolyX = Valid 0x1800000000000000000000000000c000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000000000017d
instance LFSR_Polys 150 where
  lfsrPolyX = Valid 0x20000000000001000000000000000000000000
  lfsrPolyC = Valid 0x2000000000000000000000000000000000005b
instance LFSR_Polys 151 where
  lfsrPolyX = Valid 0x48000000000000000000000000000000000000
  lfsrPolyC = Valid 0x40000000000000000000000000000000000004
instance LFSR_Polys 152 where
  lfsrPolyX = Valid 0xc0000000000000006000000000000000000000
  lfsrPolyC = Valid 0x80000000000000000000000000000000000026
instance LFSR_Polys 153 where
  lfsrPolyX = Valid 0x180000000000000000000000000000000000000
  lfsrPolyC = Valid 0x100000000000000000000000000000000000001
instance LFSR_Polys 154 where
  lfsrPolyX = Valid 0x280000000000000000000000000000005000000
  lfsrPolyC = Valid 0x200000000000000000000000000000000000076
instance LFSR_Polys 155 where
  lfsrPolyX = Valid 0x60000000c000000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000000000058
instance LFSR_Polys 156 where
  lfsrPolyX = Valid 0xc00000000000000000000000000018000000000
  lfsrPolyC = Valid 0x800000000000000000000000000000000000114
instance LFSR_Polys 157 where
  lfsrPolyX = Valid 0x1800000600000000000000000000000000000000
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000032
instance LFSR_Polys 158 where
  lfsrPolyX = Valid 0x3000000c00000000000000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000000000000009b
instance LFSR_Polys 159 where
  lfsrPolyX = Valid 0x4000000080000000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000000000003d
instance LFSR_Polys 160 where
  lfsrPolyX = Valid 0xc000300000000000000000000000000000000000
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000016
instance LFSR_Polys 161 where
  lfsrPolyX = Valid 0x10000400000000000000000000000000000000000
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000026
instance LFSR_Polys 162 where
  lfsrPolyX = Valid 0x30000000000000000000006000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000c8
instance LFSR_Polys 163 where
  lfsrPolyX = Valid 0x600000000000000c0000000000000000000000000
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000064
instance LFSR_Polys 164 where
  lfsrPolyX = Valid 0xc0060000000000000000000000000000000000000
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000f7
instance LFSR_Polys 165 where
  lfsrPolyX = Valid 0x180000006000000000000000000000000000000000
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000012d
instance LFSR_Polys 166 where
  lfsrPolyX = Valid 0x3000000000c0000000000000000000000000000000
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000206
instance LFSR_Polys 167 where
  lfsrPolyX = Valid 0x410000000000000000000000000000000000000000
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000020
instance LFSR_Polys 168 where
  lfsrPolyX = Valid 0xa00140000000000000000000000000000000000000
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000da
instance LFSR_Polys 169 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000b0
instance LFSR_Polys 170 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000c7
instance LFSR_Polys 171 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000001f
instance LFSR_Polys 172 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000040
instance LFSR_Polys 173 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000092
instance LFSR_Polys 174 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000003e
instance LFSR_Polys 175 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000020
instance LFSR_Polys 176 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000005e
instance LFSR_Polys 177 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000016
instance LFSR_Polys 178 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000c2
instance LFSR_Polys 179 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000b
instance LFSR_Polys 180 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000b6
instance LFSR_Polys 181 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000061
instance LFSR_Polys 182 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000a1
instance LFSR_Polys 183 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000c8
instance LFSR_Polys 184 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000ae
instance LFSR_Polys 185 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000085
instance LFSR_Polys 186 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000ce
instance LFSR_Polys 187 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000070
instance LFSR_Polys 188 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000032
instance LFSR_Polys 189 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000032
instance LFSR_Polys 190 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000014b
instance LFSR_Polys 191 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000005d
instance LFSR_Polys 192 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000ae
instance LFSR_Polys 193 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000fb
instance LFSR_Polys 194 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000e
instance LFSR_Polys 195 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000005b
instance LFSR_Polys 196 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000001c9
instance LFSR_Polys 197 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000f7
instance LFSR_Polys 198 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000003b9
instance LFSR_Polys 199 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000076
instance LFSR_Polys 200 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000016
instance LFSR_Polys 201 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000026
instance LFSR_Polys 202 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000068
instance LFSR_Polys 203 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000c1
instance LFSR_Polys 204 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000d5
instance LFSR_Polys 205 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000112
instance LFSR_Polys 206 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000057
instance LFSR_Polys 207 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000121
instance LFSR_Polys 208 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000e9
instance LFSR_Polys 209 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000016
instance LFSR_Polys 210 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000013a
instance LFSR_Polys 211 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000135
instance LFSR_Polys 212 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000004c
instance LFSR_Polys 213 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000032
instance LFSR_Polys 214 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000015
instance LFSR_Polys 215 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000034
instance LFSR_Polys 216 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000045
instance LFSR_Polys 217 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000038
instance LFSR_Polys 218 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000007a
instance LFSR_Polys 219 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000007a
instance LFSR_Polys 220 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000008f
instance LFSR_Polys 221 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 222 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000092
instance LFSR_Polys 223 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000001a
instance LFSR_Polys 224 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000da
instance LFSR_Polys 225 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000b6
instance LFSR_Polys 226 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 227 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 228 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 229 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000133
instance LFSR_Polys 230 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000e0
instance LFSR_Polys 231 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000004a
instance LFSR_Polys 232 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000014b
instance LFSR_Polys 233 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000005e
instance LFSR_Polys 234 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000e5
instance LFSR_Polys 235 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000e6
instance LFSR_Polys 236 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 237 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 238 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000013
instance LFSR_Polys 239 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 240 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000094
instance LFSR_Polys 241 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000bc
instance LFSR_Polys 242 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000b9
instance LFSR_Polys 243 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000091
instance LFSR_Polys 244 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 245 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000029
instance LFSR_Polys 246 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000026c
instance LFSR_Polys 247 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000010a
instance LFSR_Polys 248 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000009e
instance LFSR_Polys 249 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 250 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000037
instance LFSR_Polys 251 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000004a
instance LFSR_Polys 252 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000001b8
instance LFSR_Polys 253 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 254 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000043
instance LFSR_Polys 255 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000016
instance LFSR_Polys 256 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000212
instance LFSR_Polys 257 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000005e
instance LFSR_Polys 258 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000128
instance LFSR_Polys 259 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000fd
instance LFSR_Polys 260 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000c7
instance LFSR_Polys 261 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000068
instance LFSR_Polys 262 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000188
instance LFSR_Polys 263 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000013f
instance LFSR_Polys 264 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000301
instance LFSR_Polys 265 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000016
instance LFSR_Polys 266 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000057
instance LFSR_Polys 267 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000a4
instance LFSR_Polys 268 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000001c3
instance LFSR_Polys 269 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 270 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000ae
instance LFSR_Polys 271 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000008f
instance LFSR_Polys 272 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 273 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000043
instance LFSR_Polys 274 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 275 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 276 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000025
instance LFSR_Polys 277 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000005b
instance LFSR_Polys 278 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 279 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 280 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000112
instance LFSR_Polys 281 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000109
instance LFSR_Polys 282 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000001d4
instance LFSR_Polys 283 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 284 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000b0
instance LFSR_Polys 285 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000250
instance LFSR_Polys 286 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000fd
instance LFSR_Polys 287 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000032
instance LFSR_Polys 288 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000153
instance LFSR_Polys 289 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000007a
instance LFSR_Polys 290 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000016
instance LFSR_Polys 291 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 292 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000045
instance LFSR_Polys 293 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000012d
instance LFSR_Polys 294 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000ef
instance LFSR_Polys 295 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000001a
instance LFSR_Polys 296 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000002e1
instance LFSR_Polys 297 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 298 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 299 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000057
instance LFSR_Polys 300 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000040
instance LFSR_Polys 301 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 302 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 303 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000e3
instance LFSR_Polys 304 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 305 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000062
instance LFSR_Polys 306 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000045
instance LFSR_Polys 307 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000008a
instance LFSR_Polys 308 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000307
instance LFSR_Polys 309 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000b9
instance LFSR_Polys 310 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000091
instance LFSR_Polys 311 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000054
instance LFSR_Polys 312 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000003a8
instance LFSR_Polys 313 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000045
instance LFSR_Polys 314 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 315 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 316 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000001db
instance LFSR_Polys 317 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000004a
instance LFSR_Polys 318 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000b0
instance LFSR_Polys 319 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000097
instance LFSR_Polys 320 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000d
instance LFSR_Polys 321 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000052
instance LFSR_Polys 322 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000017b
instance LFSR_Polys 323 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 324 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000002c
instance LFSR_Polys 325 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000ab
instance LFSR_Polys 326 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000205
instance LFSR_Polys 327 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000076
instance LFSR_Polys 328 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000150
instance LFSR_Polys 329 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000009e
instance LFSR_Polys 330 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000037
instance LFSR_Polys 331 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000007a
instance LFSR_Polys 332 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000001e8
instance LFSR_Polys 333 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000002
instance LFSR_Polys 334 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 335 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000199
instance LFSR_Polys 336 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 337 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000073
instance LFSR_Polys 338 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000026
instance LFSR_Polys 339 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000057
instance LFSR_Polys 340 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000165
instance LFSR_Polys 341 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000008f
instance LFSR_Polys 342 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000ae
instance LFSR_Polys 343 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000001ed
instance LFSR_Polys 344 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000025c
instance LFSR_Polys 345 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000008a
instance LFSR_Polys 346 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000153
instance LFSR_Polys 347 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000007a
instance LFSR_Polys 348 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8
instance LFSR_Polys 349 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000032
instance LFSR_Polys 350 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000005e
instance LFSR_Polys 351 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000a4
instance LFSR_Polys 352 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000005e
instance LFSR_Polys 353 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000148
instance LFSR_Polys 354 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000195
instance LFSR_Polys 355 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000031
instance LFSR_Polys 356 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000f8
instance LFSR_Polys 357 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f8
instance LFSR_Polys 358 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b5
instance LFSR_Polys 359 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 360 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000009ad
instance LFSR_Polys 361 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 362 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000cd
instance LFSR_Polys 363 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000094
instance LFSR_Polys 364 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000028d
instance LFSR_Polys 365 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000130
instance LFSR_Polys 366 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ec
instance LFSR_Polys 367 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005d
instance LFSR_Polys 368 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 369 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002f5
instance LFSR_Polys 370 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000016
instance LFSR_Polys 371 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000086
instance LFSR_Polys 372 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b6
instance LFSR_Polys 373 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c2
instance LFSR_Polys 374 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b0
instance LFSR_Polys 375 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c1
instance LFSR_Polys 376 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d0
instance LFSR_Polys 377 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000085
instance LFSR_Polys 378 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001c3
instance LFSR_Polys 379 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000195
instance LFSR_Polys 380 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000343
instance LFSR_Polys 381 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013
instance LFSR_Polys 382 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001f6
instance LFSR_Polys 383 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111
instance LFSR_Polys 384 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022e
instance LFSR_Polys 385 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020
instance LFSR_Polys 386 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ff
instance LFSR_Polys 387 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000182
instance LFSR_Polys 388 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000019a
instance LFSR_Polys 389 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000067
instance LFSR_Polys 390 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003cb
instance LFSR_Polys 391 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000023
instance LFSR_Polys 392 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000cd
instance LFSR_Polys 393 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040
instance LFSR_Polys 394 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c2
instance LFSR_Polys 395 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fb
instance LFSR_Polys 396 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068
instance LFSR_Polys 397 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 398 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002a9
instance LFSR_Polys 399 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012b
instance LFSR_Polys 400 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000016
instance LFSR_Polys 401 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005d
instance LFSR_Polys 402 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 403 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000190
instance LFSR_Polys 404 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068
instance LFSR_Polys 405 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001aa
instance LFSR_Polys 406 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003c7
instance LFSR_Polys 407 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d3
instance LFSR_Polys 408 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002f
instance LFSR_Polys 409 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000054
instance LFSR_Polys 410 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020c
instance LFSR_Polys 411 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b6
instance LFSR_Polys 412 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ed
instance LFSR_Polys 413 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006b
instance LFSR_Polys 414 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000035b
instance LFSR_Polys 415 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010a
instance LFSR_Polys 416 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000112
instance LFSR_Polys 417 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 418 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002e8
instance LFSR_Polys 419 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013f
instance LFSR_Polys 420 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b9
instance LFSR_Polys 421 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a
instance LFSR_Polys 422 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005d
instance LFSR_Polys 423 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010f
instance LFSR_Polys 424 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d6
instance LFSR_Polys 425 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 426 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a13
instance LFSR_Polys 427 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 428 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000406
instance LFSR_Polys 429 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001c6
instance LFSR_Polys 430 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009e
instance LFSR_Polys 431 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015
instance LFSR_Polys 432 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000594
instance LFSR_Polys 433 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001b7
instance LFSR_Polys 434 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000073
instance LFSR_Polys 435 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000235
instance LFSR_Polys 436 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038
instance LFSR_Polys 437 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000023
instance LFSR_Polys 438 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000325
instance LFSR_Polys 439 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000086
instance LFSR_Polys 440 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d
instance LFSR_Polys 441 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000bc
instance LFSR_Polys 442 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000052
instance LFSR_Polys 443 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c7
instance LFSR_Polys 444 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015f
instance LFSR_Polys 445 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068
instance LFSR_Polys 446 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000351
instance LFSR_Polys 447 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ce
instance LFSR_Polys 448 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000295
instance LFSR_Polys 449 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013f
instance LFSR_Polys 450 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ea
instance LFSR_Polys 451 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000019a
instance LFSR_Polys 452 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038
instance LFSR_Polys 453 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003f8
instance LFSR_Polys 454 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011b
instance LFSR_Polys 455 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000178
instance LFSR_Polys 456 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000459
instance LFSR_Polys 457 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000136
instance LFSR_Polys 458 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010f
instance LFSR_Polys 459 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006d
instance LFSR_Polys 460 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111
instance LFSR_Polys 461 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 462 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002d2
instance LFSR_Polys 463 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002ca
instance LFSR_Polys 464 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012b
instance LFSR_Polys 465 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000086
instance LFSR_Polys 466 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e4
instance LFSR_Polys 467 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000421
instance LFSR_Polys 468 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002af
instance LFSR_Polys 469 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003e
instance LFSR_Polys 470 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009e
instance LFSR_Polys 471 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001
instance LFSR_Polys 472 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000364
instance LFSR_Polys 473 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a4
instance LFSR_Polys 474 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015c
instance LFSR_Polys 475 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000188
instance LFSR_Polys 476 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000281
instance LFSR_Polys 477 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000bc
instance LFSR_Polys 478 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000029
instance LFSR_Polys 479 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fe
instance LFSR_Polys 480 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006e
instance LFSR_Polys 481 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000014b
instance LFSR_Polys 482 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000130
instance LFSR_Polys 483 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006d
instance LFSR_Polys 484 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a9
instance LFSR_Polys 485 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d6
instance LFSR_Polys 486 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007c
instance LFSR_Polys 487 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010a
instance LFSR_Polys 488 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d
instance LFSR_Polys 489 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000130
instance LFSR_Polys 490 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000150
instance LFSR_Polys 491 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 492 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b6
instance LFSR_Polys 493 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000127
instance LFSR_Polys 494 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000379
instance LFSR_Polys 495 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030d
instance LFSR_Polys 496 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000cb
instance LFSR_Polys 497 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000351
instance LFSR_Polys 498 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fe
instance LFSR_Polys 499 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000166
instance LFSR_Polys 500 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 501 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a
instance LFSR_Polys 502 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000098
instance LFSR_Polys 503 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004
instance LFSR_Polys 504 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002f
instance LFSR_Polys 505 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018e
instance LFSR_Polys 506 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018b
instance LFSR_Polys 507 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007a
instance LFSR_Polys 508 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004f
instance LFSR_Polys 509 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c4
instance LFSR_Polys 510 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000bc
instance LFSR_Polys 511 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200
instance LFSR_Polys 512 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000092
instance LFSR_Polys 513 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 514 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000054
instance LFSR_Polys 515 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a6
instance LFSR_Polys 516 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000052
instance LFSR_Polys 517 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000316
instance LFSR_Polys 518 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001de
instance LFSR_Polys 519 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b5
instance LFSR_Polys 520 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003b6
instance LFSR_Polys 521 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000135
instance LFSR_Polys 522 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fe
instance LFSR_Polys 523 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011b
instance LFSR_Polys 524 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111
instance LFSR_Polys 525 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000029
instance LFSR_Polys 526 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111
instance LFSR_Polys 527 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000141
instance LFSR_Polys 528 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000422
instance LFSR_Polys 529 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 530 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000244
instance LFSR_Polys 531 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024b
instance LFSR_Polys 532 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001
instance LFSR_Polys 533 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e
instance LFSR_Polys 534 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000051
instance LFSR_Polys 535 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a2
instance LFSR_Polys 536 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000054
instance LFSR_Polys 537 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000203
instance LFSR_Polys 538 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013
instance LFSR_Polys 539 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000218
instance LFSR_Polys 540 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000424
instance LFSR_Polys 541 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012e
instance LFSR_Polys 542 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000106
instance LFSR_Polys 543 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038c
instance LFSR_Polys 544 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000299
instance LFSR_Polys 545 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e3
instance LFSR_Polys 546 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003b
instance LFSR_Polys 547 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f8
instance LFSR_Polys 548 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018d
instance LFSR_Polys 549 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001c3
instance LFSR_Polys 550 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ce
instance LFSR_Polys 551 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000109
instance LFSR_Polys 552 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008f9
instance LFSR_Polys 553 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003ec
instance LFSR_Polys 554 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000484
instance LFSR_Polys 555 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001fc
instance LFSR_Polys 556 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ef
instance LFSR_Polys 557 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000067
instance LFSR_Polys 558 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000272
instance LFSR_Polys 559 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000142
instance LFSR_Polys 560 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013c
instance LFSR_Polys 561 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000178
instance LFSR_Polys 562 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d6
instance LFSR_Polys 563 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d5
instance LFSR_Polys 564 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000025
instance LFSR_Polys 565 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021e
instance LFSR_Polys 566 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032
instance LFSR_Polys 567 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000036d
instance LFSR_Polys 568 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000964
instance LFSR_Polys 569 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050b
instance LFSR_Polys 570 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000073
instance LFSR_Polys 571 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000212
instance LFSR_Polys 572 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001af
instance LFSR_Polys 573 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001de
instance LFSR_Polys 574 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001dd
instance LFSR_Polys 575 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000034
instance LFSR_Polys 576 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007b7
instance LFSR_Polys 577 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000086
instance LFSR_Polys 578 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000398
instance LFSR_Polys 579 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000379
instance LFSR_Polys 580 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000029
instance LFSR_Polys 581 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002e2
instance LFSR_Polys 582 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013f
instance LFSR_Polys 583 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a2
instance LFSR_Polys 584 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d6
instance LFSR_Polys 585 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000086
instance LFSR_Polys 586 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000052
instance LFSR_Polys 587 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000421
instance LFSR_Polys 588 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003d0
instance LFSR_Polys 589 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020c
instance LFSR_Polys 590 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ad
instance LFSR_Polys 591 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000128
instance LFSR_Polys 592 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000015a
instance LFSR_Polys 593 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 594 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002af
instance LFSR_Polys 595 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000103
instance LFSR_Polys 596 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038
instance LFSR_Polys 597 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000227
instance LFSR_Polys 598 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 599 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003b
instance LFSR_Polys 600 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000601
instance LFSR_Polys 601 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004f
instance LFSR_Polys 602 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001f3
instance LFSR_Polys 603 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002c
instance LFSR_Polys 604 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000165
instance LFSR_Polys 605 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b9
instance LFSR_Polys 606 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000042b
instance LFSR_Polys 607 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000165
instance LFSR_Polys 608 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000045f
instance LFSR_Polys 609 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 610 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000043c
instance LFSR_Polys 611 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006b
instance LFSR_Polys 612 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018d
instance LFSR_Polys 613 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000022d
instance LFSR_Polys 614 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000043
instance LFSR_Polys 615 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 616 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000052f
instance LFSR_Polys 617 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ff
instance LFSR_Polys 618 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000562
instance LFSR_Polys 619 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 620 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000103
instance LFSR_Polys 621 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032c
instance LFSR_Polys 622 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001af
instance LFSR_Polys 623 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000233
instance LFSR_Polys 624 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000017b
instance LFSR_Polys 625 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000012e
instance LFSR_Polys 626 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024e
instance LFSR_Polys 627 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003e
instance LFSR_Polys 628 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002a3
instance LFSR_Polys 629 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032
instance LFSR_Polys 630 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a
instance LFSR_Polys 631 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000217
instance LFSR_Polys 632 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003d6
instance LFSR_Polys 633 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000043
instance LFSR_Polys 634 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000054
instance LFSR_Polys 635 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000fb
instance LFSR_Polys 636 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000057a
instance LFSR_Polys 637 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d5
instance LFSR_Polys 638 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000031
instance LFSR_Polys 639 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e6
instance LFSR_Polys 640 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004cf
instance LFSR_Polys 641 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ad
instance LFSR_Polys 642 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000320
instance LFSR_Polys 643 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001b7
instance LFSR_Polys 644 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005ae
instance LFSR_Polys 645 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024b
instance LFSR_Polys 646 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000166
instance LFSR_Polys 647 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 648 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000436
instance LFSR_Polys 649 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000411
instance LFSR_Polys 650 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004
instance LFSR_Polys 651 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011b
instance LFSR_Polys 652 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000076
instance LFSR_Polys 653 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f8
instance LFSR_Polys 654 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 655 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 656 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008c9
instance LFSR_Polys 657 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c1
instance LFSR_Polys 658 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000059e
instance LFSR_Polys 659 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000147
instance LFSR_Polys 660 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000080c
instance LFSR_Polys 661 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b3
instance LFSR_Polys 662 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000047b
instance LFSR_Polys 663 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002a5
instance LFSR_Polys 664 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002bb
instance LFSR_Polys 665 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000375
instance LFSR_Polys 666 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000217
instance LFSR_Polys 667 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006b3
instance LFSR_Polys 668 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000193
instance LFSR_Polys 669 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a
instance LFSR_Polys 670 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000031
instance LFSR_Polys 671 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000122
instance LFSR_Polys 672 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000037
instance LFSR_Polys 673 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ac
instance LFSR_Polys 674 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002c5
instance LFSR_Polys 675 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000025
instance LFSR_Polys 676 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024d
instance LFSR_Polys 677 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008c
instance LFSR_Polys 678 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000dc
instance LFSR_Polys 679 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 680 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e4
instance LFSR_Polys 681 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b6
instance LFSR_Polys 682 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000045
instance LFSR_Polys 683 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000018b
instance LFSR_Polys 684 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a6
instance LFSR_Polys 685 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d
instance LFSR_Polys 686 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003d9
instance LFSR_Polys 687 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000455
instance LFSR_Polys 688 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000793
instance LFSR_Polys 689 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a4
instance LFSR_Polys 690 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013a
instance LFSR_Polys 691 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ce
instance LFSR_Polys 692 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000031a
instance LFSR_Polys 693 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 694 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000256
instance LFSR_Polys 695 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000109
instance LFSR_Polys 696 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000153
instance LFSR_Polys 697 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000165
instance LFSR_Polys 698 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000033d
instance LFSR_Polys 699 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000bf
instance LFSR_Polys 700 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032
instance LFSR_Polys 701 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ca
instance LFSR_Polys 702 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000045
instance LFSR_Polys 703 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001b1
instance LFSR_Polys 704 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d6
instance LFSR_Polys 705 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b0
instance LFSR_Polys 706 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021d
instance LFSR_Polys 707 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e8
instance LFSR_Polys 708 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a
instance LFSR_Polys 709 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d
instance LFSR_Polys 710 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003cb
instance LFSR_Polys 711 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002f0
instance LFSR_Polys 712 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001c
instance LFSR_Polys 713 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000534
instance LFSR_Polys 714 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004fc
instance LFSR_Polys 715 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000049
instance LFSR_Polys 716 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000472
instance LFSR_Polys 717 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000573
instance LFSR_Polys 718 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013
instance LFSR_Polys 719 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000029f
instance LFSR_Polys 720 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000482
instance LFSR_Polys 721 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000bc
instance LFSR_Polys 722 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003b
instance LFSR_Polys 723 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001c6
instance LFSR_Polys 724 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006f2
instance LFSR_Polys 725 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d5
instance LFSR_Polys 726 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 727 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000195
instance LFSR_Polys 728 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e
instance LFSR_Polys 729 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000136
instance LFSR_Polys 730 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b2d
instance LFSR_Polys 731 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 732 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004c
instance LFSR_Polys 733 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c2
instance LFSR_Polys 734 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004a9
instance LFSR_Polys 735 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c2
instance LFSR_Polys 736 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000493
instance LFSR_Polys 737 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010
instance LFSR_Polys 738 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000178
instance LFSR_Polys 739 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001d2
instance LFSR_Polys 740 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000319
instance LFSR_Polys 741 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000184
instance LFSR_Polys 742 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000570
instance LFSR_Polys 743 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000379
instance LFSR_Polys 744 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011b
instance LFSR_Polys 745 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d0
instance LFSR_Polys 746 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000057
instance LFSR_Polys 747 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000228
instance LFSR_Polys 748 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006c7
instance LFSR_Polys 749 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 750 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003e3
instance LFSR_Polys 751 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000079
instance LFSR_Polys 752 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000023a
instance LFSR_Polys 753 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000172
instance LFSR_Polys 754 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000925
instance LFSR_Polys 755 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006df
instance LFSR_Polys 756 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000090b
instance LFSR_Polys 757 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 758 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007a3
instance LFSR_Polys 759 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000106
instance LFSR_Polys 760 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000067c
instance LFSR_Polys 761 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004
instance LFSR_Polys 762 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 763 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 764 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000034
instance LFSR_Polys 765 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002d8
instance LFSR_Polys 766 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005bf
instance LFSR_Polys 767 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8
instance LFSR_Polys 768 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010d4
instance LFSR_Polys 769 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000160
instance LFSR_Polys 770 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000070a
instance LFSR_Polys 771 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a9
instance LFSR_Polys 772 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040
instance LFSR_Polys 773 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002a0
instance LFSR_Polys 774 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a7
instance LFSR_Polys 775 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068
instance LFSR_Polys 776 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000664
instance LFSR_Polys 777 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000398
instance LFSR_Polys 778 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ea
instance LFSR_Polys 779 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000227
instance LFSR_Polys 780 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000ef
instance LFSR_Polys 781 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000236
instance LFSR_Polys 782 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006b
instance LFSR_Polys 783 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001dd
instance LFSR_Polys 784 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000048e
instance LFSR_Polys 785 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005e
instance LFSR_Polys 786 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002b4
instance LFSR_Polys 787 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000064
instance LFSR_Polys 788 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003e5
instance LFSR_Polys 789 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013
instance LFSR_Polys 790 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000144
instance LFSR_Polys 791 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000029
instance LFSR_Polys 792 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000139
instance LFSR_Polys 793 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000109
instance LFSR_Polys 794 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000023c
instance LFSR_Polys 795 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030e
instance LFSR_Polys 796 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f1
instance LFSR_Polys 797 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002aa
instance LFSR_Polys 798 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000064
instance LFSR_Polys 799 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000bc
instance LFSR_Polys 800 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000166
instance LFSR_Polys 801 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000141
instance LFSR_Polys 802 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ed
instance LFSR_Polys 803 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d5
instance LFSR_Polys 804 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000340
instance LFSR_Polys 805 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000076
instance LFSR_Polys 806 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000310
instance LFSR_Polys 807 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000040
instance LFSR_Polys 808 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ed
instance LFSR_Polys 809 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000085
instance LFSR_Polys 810 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000169
instance LFSR_Polys 811 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000073
instance LFSR_Polys 812 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000077d
instance LFSR_Polys 813 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d3
instance LFSR_Polys 814 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000209
instance LFSR_Polys 815 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001ed
instance LFSR_Polys 816 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c5e
instance LFSR_Polys 817 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000287
instance LFSR_Polys 818 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000f2
instance LFSR_Polys 819 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011e
instance LFSR_Polys 820 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001af
instance LFSR_Polys 821 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000259
instance LFSR_Polys 822 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006bc
instance LFSR_Polys 823 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100
instance LFSR_Polys 824 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001f
instance LFSR_Polys 825 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003b0
instance LFSR_Polys 826 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013a
instance LFSR_Polys 827 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003d
instance LFSR_Polys 828 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030d
instance LFSR_Polys 829 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000d
instance LFSR_Polys 830 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e3
instance LFSR_Polys 831 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000153
instance LFSR_Polys 832 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e6
instance LFSR_Polys 833 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007c
instance LFSR_Polys 834 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000026f
instance LFSR_Polys 835 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002b2
instance LFSR_Polys 836 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000302
instance LFSR_Polys 837 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b0
instance LFSR_Polys 838 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000263
instance LFSR_Polys 839 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e4
instance LFSR_Polys 840 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000411
instance LFSR_Polys 841 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038
instance LFSR_Polys 842 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 843 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000033b
instance LFSR_Polys 844 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001f5
instance LFSR_Polys 845 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002
instance LFSR_Polys 846 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006d3
instance LFSR_Polys 847 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000272
instance LFSR_Polys 848 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 849 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000133
instance LFSR_Polys 850 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000697
instance LFSR_Polys 851 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000178
instance LFSR_Polys 852 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000098
instance LFSR_Polys 853 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000241
instance LFSR_Polys 854 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000054
instance LFSR_Polys 855 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000024b
instance LFSR_Polys 856 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068c
instance LFSR_Polys 857 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000034
instance LFSR_Polys 858 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004e7
instance LFSR_Polys 859 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000135
instance LFSR_Polys 860 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000199
instance LFSR_Polys 861 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000112
instance LFSR_Polys 862 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000061
instance LFSR_Polys 863 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000026
instance LFSR_Polys 864 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001b52
instance LFSR_Polys 865 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001
instance LFSR_Polys 866 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000263
instance LFSR_Polys 867 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000112
instance LFSR_Polys 868 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000050e
instance LFSR_Polys 869 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000036e
instance LFSR_Polys 870 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000081b
instance LFSR_Polys 871 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000239
instance LFSR_Polys 872 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002ed
instance LFSR_Polys 873 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000045
instance LFSR_Polys 874 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000781
instance LFSR_Polys 875 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007d8
instance LFSR_Polys 876 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000871
instance LFSR_Polys 877 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000038
instance LFSR_Polys 878 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002b1
instance LFSR_Polys 879 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000114
instance LFSR_Polys 880 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000546
instance LFSR_Polys 881 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000490
instance LFSR_Polys 882 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000411
instance LFSR_Polys 883 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001a3
instance LFSR_Polys 884 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000dc
instance LFSR_Polys 885 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c1
instance LFSR_Polys 886 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000032f
instance LFSR_Polys 887 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000068
instance LFSR_Polys 888 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e7
instance LFSR_Polys 889 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001dd
instance LFSR_Polys 890 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000054c
instance LFSR_Polys 891 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000da
instance LFSR_Polys 892 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000439
instance LFSR_Polys 893 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 894 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009b
instance LFSR_Polys 895 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009d
instance LFSR_Polys 896 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000295
instance LFSR_Polys 897 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000039d
instance LFSR_Polys 898 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002cf
instance LFSR_Polys 899 where
  lfsrPolyC = Valid 0x400000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000439
instance LFSR_Polys 900 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001
instance LFSR_Polys 901 where
  lfsrPolyC = Valid 0x1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000357
instance LFSR_Polys 902 where
  lfsrPolyC = Valid 0x20000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000e3
instance LFSR_Polys 903 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c1
instance LFSR_Polys 904 where
  lfsrPolyC = Valid 0x8000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000711
instance LFSR_Polys 905 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000135
instance LFSR_Polys 906 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000004b4
instance LFSR_Polys 907 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000017d
instance LFSR_Polys 908 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000c8
instance LFSR_Polys 909 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000373
instance LFSR_Polys 910 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005c8
instance LFSR_Polys 911 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a1
instance LFSR_Polys 912 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000baf
instance LFSR_Polys 913 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000030d
instance LFSR_Polys 914 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000b
instance LFSR_Polys 915 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000a4
instance LFSR_Polys 916 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000031a
instance LFSR_Polys 917 where
  lfsrPolyC = Valid 0x100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000005c8
instance LFSR_Polys 918 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000003c7
instance LFSR_Polys 919 where
  lfsrPolyC = Valid 0x40000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000150
instance LFSR_Polys 920 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000469
instance LFSR_Polys 921 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000013a
instance LFSR_Polys 922 where
  lfsrPolyC = Valid 0x200000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000070
instance LFSR_Polys 923 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001e1
instance LFSR_Polys 924 where
  lfsrPolyC = Valid 0x800000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000592
instance LFSR_Polys 925 where
  lfsrPolyC = Valid 0x10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000df
instance LFSR_Polys 926 where
  lfsrPolyC = Valid 0x2000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000525
instance LFSR_Polys 927 where
  lfsrPolyC = Valid 0x4000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000144
instance LFSR_Polys 928 where
  lfsrPolyC = Valid 0x80000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007d8

-- Define functions similar to those in LFSR.bs for backward compatibility. The
-- entries for 4, 8, 16, and 32 are already defined in LFSR.bs (with the same K
-- polynomials), but they are defined here anyway for completeness.

-- TODO: Do we even want these? I don't think they are used, or likely to be.

mkLFSR_2 :: (IsModule m c) => m (LFSR (Bit 2))
mkLFSR_2 = mkLFSR
mkLFSR_3 :: (IsModule m c) => m (LFSR (Bit 3))
mkLFSR_3 = mkLFSR
mkLFSR_4 :: (IsModule m c) => m (LFSR (Bit 4))
mkLFSR_4 = mkLFSR
mkLFSR_5 :: (IsModule m c) => m (LFSR (Bit 5))
mkLFSR_5 = mkLFSR
mkLFSR_6 :: (IsModule m c) => m (LFSR (Bit 6))
mkLFSR_6 = mkLFSR
mkLFSR_7 :: (IsModule m c) => m (LFSR (Bit 7))
mkLFSR_7 = mkLFSR
mkLFSR_8 :: (IsModule m c) => m (LFSR (Bit 8))
mkLFSR_8 = mkLFSR
mkLFSR_9 :: (IsModule m c) => m (LFSR (Bit 9))
mkLFSR_9 = mkLFSR
mkLFSR_10 :: (IsModule m c) => m (LFSR (Bit 10))
mkLFSR_10 = mkLFSR
mkLFSR_11 :: (IsModule m c) => m (LFSR (Bit 11))
mkLFSR_11 = mkLFSR
mkLFSR_12 :: (IsModule m c) => m (LFSR (Bit 12))
mkLFSR_12 = mkLFSR
mkLFSR_13 :: (IsModule m c) => m (LFSR (Bit 13))
mkLFSR_13 = mkLFSR
mkLFSR_14 :: (IsModule m c) => m (LFSR (Bit 14))
mkLFSR_14 = mkLFSR
mkLFSR_15 :: (IsModule m c) => m (LFSR (Bit 15))
mkLFSR_15 = mkLFSR
mkLFSR_16 :: (IsModule m c) => m (LFSR (Bit 16))
mkLFSR_16 = mkLFSR
mkLFSR_17 :: (IsModule m c) => m (LFSR (Bit 17))
mkLFSR_17 = mkLFSR
mkLFSR_18 :: (IsModule m c) => m (LFSR (Bit 18))
mkLFSR_18 = mkLFSR
mkLFSR_19 :: (IsModule m c) => m (LFSR (Bit 19))
mkLFSR_19 = mkLFSR
mkLFSR_20 :: (IsModule m c) => m (LFSR (Bit 20))
mkLFSR_20 = mkLFSR
mkLFSR_21 :: (IsModule m c) => m (LFSR (Bit 21))
mkLFSR_21 = mkLFSR
mkLFSR_22 :: (IsModule m c) => m (LFSR (Bit 22))
mkLFSR_22 = mkLFSR
mkLFSR_23 :: (IsModule m c) => m (LFSR (Bit 23))
mkLFSR_23 = mkLFSR
mkLFSR_24 :: (IsModule m c) => m (LFSR (Bit 24))
mkLFSR_24 = mkLFSR
mkLFSR_25 :: (IsModule m c) => m (LFSR (Bit 25))
mkLFSR_25 = mkLFSR
mkLFSR_26 :: (IsModule m c) => m (LFSR (Bit 26))
mkLFSR_26 = mkLFSR
mkLFSR_27 :: (IsModule m c) => m (LFSR (Bit 27))
mkLFSR_27 = mkLFSR
mkLFSR_28 :: (IsModule m c) => m (LFSR (Bit 28))
mkLFSR_28 = mkLFSR
mkLFSR_29 :: (IsModule m c) => m (LFSR (Bit 29))
mkLFSR_29 = mkLFSR
mkLFSR_30 :: (IsModule m c) => m (LFSR (Bit 30))
mkLFSR_30 = mkLFSR
mkLFSR_31 :: (IsModule m c) => m (LFSR (Bit 31))
mkLFSR_31 = mkLFSR
mkLFSR_32 :: (IsModule m c) => m (LFSR (Bit 32))
mkLFSR_32 = mkLFSR
mkLFSR_33 :: (IsModule m c) => m (LFSR (Bit 33))
mkLFSR_33 = mkLFSR
mkLFSR_34 :: (IsModule m c) => m (LFSR (Bit 34))
mkLFSR_34 = mkLFSR
mkLFSR_35 :: (IsModule m c) => m (LFSR (Bit 35))
mkLFSR_35 = mkLFSR
mkLFSR_36 :: (IsModule m c) => m (LFSR (Bit 36))
mkLFSR_36 = mkLFSR
mkLFSR_37 :: (IsModule m c) => m (LFSR (Bit 37))
mkLFSR_37 = mkLFSR
mkLFSR_38 :: (IsModule m c) => m (LFSR (Bit 38))
mkLFSR_38 = mkLFSR
mkLFSR_39 :: (IsModule m c) => m (LFSR (Bit 39))
mkLFSR_39 = mkLFSR
mkLFSR_40 :: (IsModule m c) => m (LFSR (Bit 40))
mkLFSR_40 = mkLFSR
mkLFSR_41 :: (IsModule m c) => m (LFSR (Bit 41))
mkLFSR_41 = mkLFSR
mkLFSR_42 :: (IsModule m c) => m (LFSR (Bit 42))
mkLFSR_42 = mkLFSR
mkLFSR_43 :: (IsModule m c) => m (LFSR (Bit 43))
mkLFSR_43 = mkLFSR
mkLFSR_44 :: (IsModule m c) => m (LFSR (Bit 44))
mkLFSR_44 = mkLFSR
mkLFSR_45 :: (IsModule m c) => m (LFSR (Bit 45))
mkLFSR_45 = mkLFSR
mkLFSR_46 :: (IsModule m c) => m (LFSR (Bit 46))
mkLFSR_46 = mkLFSR
mkLFSR_47 :: (IsModule m c) => m (LFSR (Bit 47))
mkLFSR_47 = mkLFSR
mkLFSR_48 :: (IsModule m c) => m (LFSR (Bit 48))
mkLFSR_48 = mkLFSR
mkLFSR_49 :: (IsModule m c) => m (LFSR (Bit 49))
mkLFSR_49 = mkLFSR
mkLFSR_50 :: (IsModule m c) => m (LFSR (Bit 50))
mkLFSR_50 = mkLFSR
mkLFSR_51 :: (IsModule m c) => m (LFSR (Bit 51))
mkLFSR_51 = mkLFSR
mkLFSR_52 :: (IsModule m c) => m (LFSR (Bit 52))
mkLFSR_52 = mkLFSR
mkLFSR_53 :: (IsModule m c) => m (LFSR (Bit 53))
mkLFSR_53 = mkLFSR
mkLFSR_54 :: (IsModule m c) => m (LFSR (Bit 54))
mkLFSR_54 = mkLFSR
mkLFSR_55 :: (IsModule m c) => m (LFSR (Bit 55))
mkLFSR_55 = mkLFSR
mkLFSR_56 :: (IsModule m c) => m (LFSR (Bit 56))
mkLFSR_56 = mkLFSR
mkLFSR_57 :: (IsModule m c) => m (LFSR (Bit 57))
mkLFSR_57 = mkLFSR
mkLFSR_58 :: (IsModule m c) => m (LFSR (Bit 58))
mkLFSR_58 = mkLFSR
mkLFSR_59 :: (IsModule m c) => m (LFSR (Bit 59))
mkLFSR_59 = mkLFSR
mkLFSR_60 :: (IsModule m c) => m (LFSR (Bit 60))
mkLFSR_60 = mkLFSR
mkLFSR_61 :: (IsModule m c) => m (LFSR (Bit 61))
mkLFSR_61 = mkLFSR
mkLFSR_62 :: (IsModule m c) => m (LFSR (Bit 62))
mkLFSR_62 = mkLFSR
mkLFSR_63 :: (IsModule m c) => m (LFSR (Bit 63))
mkLFSR_63 = mkLFSR
mkLFSR_64 :: (IsModule m c) => m (LFSR (Bit 64))
mkLFSR_64 = mkLFSR
mkLFSR_65 :: (IsModule m c) => m (LFSR (Bit 65))
mkLFSR_65 = mkLFSR
mkLFSR_66 :: (IsModule m c) => m (LFSR (Bit 66))
mkLFSR_66 = mkLFSR
mkLFSR_67 :: (IsModule m c) => m (LFSR (Bit 67))
mkLFSR_67 = mkLFSR
mkLFSR_68 :: (IsModule m c) => m (LFSR (Bit 68))
mkLFSR_68 = mkLFSR
mkLFSR_69 :: (IsModule m c) => m (LFSR (Bit 69))
mkLFSR_69 = mkLFSR
mkLFSR_70 :: (IsModule m c) => m (LFSR (Bit 70))
mkLFSR_70 = mkLFSR
mkLFSR_71 :: (IsModule m c) => m (LFSR (Bit 71))
mkLFSR_71 = mkLFSR
mkLFSR_72 :: (IsModule m c) => m (LFSR (Bit 72))
mkLFSR_72 = mkLFSR
mkLFSR_73 :: (IsModule m c) => m (LFSR (Bit 73))
mkLFSR_73 = mkLFSR
mkLFSR_74 :: (IsModule m c) => m (LFSR (Bit 74))
mkLFSR_74 = mkLFSR
mkLFSR_75 :: (IsModule m c) => m (LFSR (Bit 75))
mkLFSR_75 = mkLFSR
mkLFSR_76 :: (IsModule m c) => m (LFSR (Bit 76))
mkLFSR_76 = mkLFSR
mkLFSR_77 :: (IsModule m c) => m (LFSR (Bit 77))
mkLFSR_77 = mkLFSR
mkLFSR_78 :: (IsModule m c) => m (LFSR (Bit 78))
mkLFSR_78 = mkLFSR
mkLFSR_79 :: (IsModule m c) => m (LFSR (Bit 79))
mkLFSR_79 = mkLFSR
mkLFSR_80 :: (IsModule m c) => m (LFSR (Bit 80))
mkLFSR_80 = mkLFSR
mkLFSR_81 :: (IsModule m c) => m (LFSR (Bit 81))
mkLFSR_81 = mkLFSR
mkLFSR_82 :: (IsModule m c) => m (LFSR (Bit 82))
mkLFSR_82 = mkLFSR
mkLFSR_83 :: (IsModule m c) => m (LFSR (Bit 83))
mkLFSR_83 = mkLFSR
mkLFSR_84 :: (IsModule m c) => m (LFSR (Bit 84))
mkLFSR_84 = mkLFSR
mkLFSR_85 :: (IsModule m c) => m (LFSR (Bit 85))
mkLFSR_85 = mkLFSR
mkLFSR_86 :: (IsModule m c) => m (LFSR (Bit 86))
mkLFSR_86 = mkLFSR
mkLFSR_87 :: (IsModule m c) => m (LFSR (Bit 87))
mkLFSR_87 = mkLFSR
mkLFSR_88 :: (IsModule m c) => m (LFSR (Bit 88))
mkLFSR_88 = mkLFSR
mkLFSR_89 :: (IsModule m c) => m (LFSR (Bit 89))
mkLFSR_89 = mkLFSR
mkLFSR_90 :: (IsModule m c) => m (LFSR (Bit 90))
mkLFSR_90 = mkLFSR
mkLFSR_91 :: (IsModule m c) => m (LFSR (Bit 91))
mkLFSR_91 = mkLFSR
mkLFSR_92 :: (IsModule m c) => m (LFSR (Bit 92))
mkLFSR_92 = mkLFSR
mkLFSR_93 :: (IsModule m c) => m (LFSR (Bit 93))
mkLFSR_93 = mkLFSR
mkLFSR_94 :: (IsModule m c) => m (LFSR (Bit 94))
mkLFSR_94 = mkLFSR
mkLFSR_95 :: (IsModule m c) => m (LFSR (Bit 95))
mkLFSR_95 = mkLFSR
mkLFSR_96 :: (IsModule m c) => m (LFSR (Bit 96))
mkLFSR_96 = mkLFSR
mkLFSR_97 :: (IsModule m c) => m (LFSR (Bit 97))
mkLFSR_97 = mkLFSR
mkLFSR_98 :: (IsModule m c) => m (LFSR (Bit 98))
mkLFSR_98 = mkLFSR
mkLFSR_99 :: (IsModule m c) => m (LFSR (Bit 99))
mkLFSR_99 = mkLFSR
mkLFSR_100 :: (IsModule m c) => m (LFSR (Bit 100))
mkLFSR_100 = mkLFSR
mkLFSR_101 :: (IsModule m c) => m (LFSR (Bit 101))
mkLFSR_101 = mkLFSR
mkLFSR_102 :: (IsModule m c) => m (LFSR (Bit 102))
mkLFSR_102 = mkLFSR
mkLFSR_103 :: (IsModule m c) => m (LFSR (Bit 103))
mkLFSR_103 = mkLFSR
mkLFSR_104 :: (IsModule m c) => m (LFSR (Bit 104))
mkLFSR_104 = mkLFSR
mkLFSR_105 :: (IsModule m c) => m (LFSR (Bit 105))
mkLFSR_105 = mkLFSR
mkLFSR_106 :: (IsModule m c) => m (LFSR (Bit 106))
mkLFSR_106 = mkLFSR
mkLFSR_107 :: (IsModule m c) => m (LFSR (Bit 107))
mkLFSR_107 = mkLFSR
mkLFSR_108 :: (IsModule m c) => m (LFSR (Bit 108))
mkLFSR_108 = mkLFSR
mkLFSR_109 :: (IsModule m c) => m (LFSR (Bit 109))
mkLFSR_109 = mkLFSR
mkLFSR_110 :: (IsModule m c) => m (LFSR (Bit 110))
mkLFSR_110 = mkLFSR
mkLFSR_111 :: (IsModule m c) => m (LFSR (Bit 111))
mkLFSR_111 = mkLFSR
mkLFSR_112 :: (IsModule m c) => m (LFSR (Bit 112))
mkLFSR_112 = mkLFSR
mkLFSR_113 :: (IsModule m c) => m (LFSR (Bit 113))
mkLFSR_113 = mkLFSR
mkLFSR_114 :: (IsModule m c) => m (LFSR (Bit 114))
mkLFSR_114 = mkLFSR
mkLFSR_115 :: (IsModule m c) => m (LFSR (Bit 115))
mkLFSR_115 = mkLFSR
mkLFSR_116 :: (IsModule m c) => m (LFSR (Bit 116))
mkLFSR_116 = mkLFSR
mkLFSR_117 :: (IsModule m c) => m (LFSR (Bit 117))
mkLFSR_117 = mkLFSR
mkLFSR_118 :: (IsModule m c) => m (LFSR (Bit 118))
mkLFSR_118 = mkLFSR
mkLFSR_119 :: (IsModule m c) => m (LFSR (Bit 119))
mkLFSR_119 = mkLFSR
mkLFSR_120 :: (IsModule m c) => m (LFSR (Bit 120))
mkLFSR_120 = mkLFSR
mkLFSR_121 :: (IsModule m c) => m (LFSR (Bit 121))
mkLFSR_121 = mkLFSR
mkLFSR_122 :: (IsModule m c) => m (LFSR (Bit 122))
mkLFSR_122 = mkLFSR
mkLFSR_123 :: (IsModule m c) => m (LFSR (Bit 123))
mkLFSR_123 = mkLFSR
mkLFSR_124 :: (IsModule m c) => m (LFSR (Bit 124))
mkLFSR_124 = mkLFSR
mkLFSR_125 :: (IsModule m c) => m (LFSR (Bit 125))
mkLFSR_125 = mkLFSR
mkLFSR_126 :: (IsModule m c) => m (LFSR (Bit 126))
mkLFSR_126 = mkLFSR
mkLFSR_127 :: (IsModule m c) => m (LFSR (Bit 127))
mkLFSR_127 = mkLFSR
mkLFSR_128 :: (IsModule m c) => m (LFSR (Bit 128))
mkLFSR_128 = mkLFSR
mkLFSR_129 :: (IsModule m c) => m (LFSR (Bit 129))
mkLFSR_129 = mkLFSR
mkLFSR_130 :: (IsModule m c) => m (LFSR (Bit 130))
mkLFSR_130 = mkLFSR
mkLFSR_131 :: (IsModule m c) => m (LFSR (Bit 131))
mkLFSR_131 = mkLFSR
mkLFSR_132 :: (IsModule m c) => m (LFSR (Bit 132))
mkLFSR_132 = mkLFSR
mkLFSR_133 :: (IsModule m c) => m (LFSR (Bit 133))
mkLFSR_133 = mkLFSR
mkLFSR_134 :: (IsModule m c) => m (LFSR (Bit 134))
mkLFSR_134 = mkLFSR
mkLFSR_135 :: (IsModule m c) => m (LFSR (Bit 135))
mkLFSR_135 = mkLFSR
mkLFSR_136 :: (IsModule m c) => m (LFSR (Bit 136))
mkLFSR_136 = mkLFSR
mkLFSR_137 :: (IsModule m c) => m (LFSR (Bit 137))
mkLFSR_137 = mkLFSR
mkLFSR_138 :: (IsModule m c) => m (LFSR (Bit 138))
mkLFSR_138 = mkLFSR
mkLFSR_139 :: (IsModule m c) => m (LFSR (Bit 139))
mkLFSR_139 = mkLFSR
mkLFSR_140 :: (IsModule m c) => m (LFSR (Bit 140))
mkLFSR_140 = mkLFSR
mkLFSR_141 :: (IsModule m c) => m (LFSR (Bit 141))
mkLFSR_141 = mkLFSR
mkLFSR_142 :: (IsModule m c) => m (LFSR (Bit 142))
mkLFSR_142 = mkLFSR
mkLFSR_143 :: (IsModule m c) => m (LFSR (Bit 143))
mkLFSR_143 = mkLFSR
mkLFSR_144 :: (IsModule m c) => m (LFSR (Bit 144))
mkLFSR_144 = mkLFSR
mkLFSR_145 :: (IsModule m c) => m (LFSR (Bit 145))
mkLFSR_145 = mkLFSR
mkLFSR_146 :: (IsModule m c) => m (LFSR (Bit 146))
mkLFSR_146 = mkLFSR
mkLFSR_147 :: (IsModule m c) => m (LFSR (Bit 147))
mkLFSR_147 = mkLFSR
mkLFSR_148 :: (IsModule m c) => m (LFSR (Bit 148))
mkLFSR_148 = mkLFSR
mkLFSR_149 :: (IsModule m c) => m (LFSR (Bit 149))
mkLFSR_149 = mkLFSR
mkLFSR_150 :: (IsModule m c) => m (LFSR (Bit 150))
mkLFSR_150 = mkLFSR
mkLFSR_151 :: (IsModule m c) => m (LFSR (Bit 151))
mkLFSR_151 = mkLFSR
mkLFSR_152 :: (IsModule m c) => m (LFSR (Bit 152))
mkLFSR_152 = mkLFSR
mkLFSR_153 :: (IsModule m c) => m (LFSR (Bit 153))
mkLFSR_153 = mkLFSR
mkLFSR_154 :: (IsModule m c) => m (LFSR (Bit 154))
mkLFSR_154 = mkLFSR
mkLFSR_155 :: (IsModule m c) => m (LFSR (Bit 155))
mkLFSR_155 = mkLFSR
mkLFSR_156 :: (IsModule m c) => m (LFSR (Bit 156))
mkLFSR_156 = mkLFSR
mkLFSR_157 :: (IsModule m c) => m (LFSR (Bit 157))
mkLFSR_157 = mkLFSR
mkLFSR_158 :: (IsModule m c) => m (LFSR (Bit 158))
mkLFSR_158 = mkLFSR
mkLFSR_159 :: (IsModule m c) => m (LFSR (Bit 159))
mkLFSR_159 = mkLFSR
mkLFSR_160 :: (IsModule m c) => m (LFSR (Bit 160))
mkLFSR_160 = mkLFSR
mkLFSR_161 :: (IsModule m c) => m (LFSR (Bit 161))
mkLFSR_161 = mkLFSR
mkLFSR_162 :: (IsModule m c) => m (LFSR (Bit 162))
mkLFSR_162 = mkLFSR
mkLFSR_163 :: (IsModule m c) => m (LFSR (Bit 163))
mkLFSR_163 = mkLFSR
mkLFSR_164 :: (IsModule m c) => m (LFSR (Bit 164))
mkLFSR_164 = mkLFSR
mkLFSR_165 :: (IsModule m c) => m (LFSR (Bit 165))
mkLFSR_165 = mkLFSR
mkLFSR_166 :: (IsModule m c) => m (LFSR (Bit 166))
mkLFSR_166 = mkLFSR
mkLFSR_167 :: (IsModule m c) => m (LFSR (Bit 167))
mkLFSR_167 = mkLFSR
mkLFSR_168 :: (IsModule m c) => m (LFSR (Bit 168))
mkLFSR_168 = mkLFSR
mkLFSR_169 :: (IsModule m c) => m (LFSR (Bit 169))
mkLFSR_169 = mkLFSR
mkLFSR_170 :: (IsModule m c) => m (LFSR (Bit 170))
mkLFSR_170 = mkLFSR
mkLFSR_171 :: (IsModule m c) => m (LFSR (Bit 171))
mkLFSR_171 = mkLFSR
mkLFSR_172 :: (IsModule m c) => m (LFSR (Bit 172))
mkLFSR_172 = mkLFSR
mkLFSR_173 :: (IsModule m c) => m (LFSR (Bit 173))
mkLFSR_173 = mkLFSR
mkLFSR_174 :: (IsModule m c) => m (LFSR (Bit 174))
mkLFSR_174 = mkLFSR
mkLFSR_175 :: (IsModule m c) => m (LFSR (Bit 175))
mkLFSR_175 = mkLFSR
mkLFSR_176 :: (IsModule m c) => m (LFSR (Bit 176))
mkLFSR_176 = mkLFSR
mkLFSR_177 :: (IsModule m c) => m (LFSR (Bit 177))
mkLFSR_177 = mkLFSR
mkLFSR_178 :: (IsModule m c) => m (LFSR (Bit 178))
mkLFSR_178 = mkLFSR
mkLFSR_179 :: (IsModule m c) => m (LFSR (Bit 179))
mkLFSR_179 = mkLFSR
mkLFSR_180 :: (IsModule m c) => m (LFSR (Bit 180))
mkLFSR_180 = mkLFSR
mkLFSR_181 :: (IsModule m c) => m (LFSR (Bit 181))
mkLFSR_181 = mkLFSR
mkLFSR_182 :: (IsModule m c) => m (LFSR (Bit 182))
mkLFSR_182 = mkLFSR
mkLFSR_183 :: (IsModule m c) => m (LFSR (Bit 183))
mkLFSR_183 = mkLFSR
mkLFSR_184 :: (IsModule m c) => m (LFSR (Bit 184))
mkLFSR_184 = mkLFSR
mkLFSR_185 :: (IsModule m c) => m (LFSR (Bit 185))
mkLFSR_185 = mkLFSR
mkLFSR_186 :: (IsModule m c) => m (LFSR (Bit 186))
mkLFSR_186 = mkLFSR
mkLFSR_187 :: (IsModule m c) => m (LFSR (Bit 187))
mkLFSR_187 = mkLFSR
mkLFSR_188 :: (IsModule m c) => m (LFSR (Bit 188))
mkLFSR_188 = mkLFSR
mkLFSR_189 :: (IsModule m c) => m (LFSR (Bit 189))
mkLFSR_189 = mkLFSR
mkLFSR_190 :: (IsModule m c) => m (LFSR (Bit 190))
mkLFSR_190 = mkLFSR
mkLFSR_191 :: (IsModule m c) => m (LFSR (Bit 191))
mkLFSR_191 = mkLFSR
mkLFSR_192 :: (IsModule m c) => m (LFSR (Bit 192))
mkLFSR_192 = mkLFSR
mkLFSR_193 :: (IsModule m c) => m (LFSR (Bit 193))
mkLFSR_193 = mkLFSR
mkLFSR_194 :: (IsModule m c) => m (LFSR (Bit 194))
mkLFSR_194 = mkLFSR
mkLFSR_195 :: (IsModule m c) => m (LFSR (Bit 195))
mkLFSR_195 = mkLFSR
mkLFSR_196 :: (IsModule m c) => m (LFSR (Bit 196))
mkLFSR_196 = mkLFSR
mkLFSR_197 :: (IsModule m c) => m (LFSR (Bit 197))
mkLFSR_197 = mkLFSR
mkLFSR_198 :: (IsModule m c) => m (LFSR (Bit 198))
mkLFSR_198 = mkLFSR
mkLFSR_199 :: (IsModule m c) => m (LFSR (Bit 199))
mkLFSR_199 = mkLFSR
mkLFSR_200 :: (IsModule m c) => m (LFSR (Bit 200))
mkLFSR_200 = mkLFSR
mkLFSR_201 :: (IsModule m c) => m (LFSR (Bit 201))
mkLFSR_201 = mkLFSR
mkLFSR_202 :: (IsModule m c) => m (LFSR (Bit 202))
mkLFSR_202 = mkLFSR
mkLFSR_203 :: (IsModule m c) => m (LFSR (Bit 203))
mkLFSR_203 = mkLFSR
mkLFSR_204 :: (IsModule m c) => m (LFSR (Bit 204))
mkLFSR_204 = mkLFSR
mkLFSR_205 :: (IsModule m c) => m (LFSR (Bit 205))
mkLFSR_205 = mkLFSR
mkLFSR_206 :: (IsModule m c) => m (LFSR (Bit 206))
mkLFSR_206 = mkLFSR
mkLFSR_207 :: (IsModule m c) => m (LFSR (Bit 207))
mkLFSR_207 = mkLFSR
mkLFSR_208 :: (IsModule m c) => m (LFSR (Bit 208))
mkLFSR_208 = mkLFSR
mkLFSR_209 :: (IsModule m c) => m (LFSR (Bit 209))
mkLFSR_209 = mkLFSR
mkLFSR_210 :: (IsModule m c) => m (LFSR (Bit 210))
mkLFSR_210 = mkLFSR
mkLFSR_211 :: (IsModule m c) => m (LFSR (Bit 211))
mkLFSR_211 = mkLFSR
mkLFSR_212 :: (IsModule m c) => m (LFSR (Bit 212))
mkLFSR_212 = mkLFSR
mkLFSR_213 :: (IsModule m c) => m (LFSR (Bit 213))
mkLFSR_213 = mkLFSR
mkLFSR_214 :: (IsModule m c) => m (LFSR (Bit 214))
mkLFSR_214 = mkLFSR
mkLFSR_215 :: (IsModule m c) => m (LFSR (Bit 215))
mkLFSR_215 = mkLFSR
mkLFSR_216 :: (IsModule m c) => m (LFSR (Bit 216))
mkLFSR_216 = mkLFSR
mkLFSR_217 :: (IsModule m c) => m (LFSR (Bit 217))
mkLFSR_217 = mkLFSR
mkLFSR_218 :: (IsModule m c) => m (LFSR (Bit 218))
mkLFSR_218 = mkLFSR
mkLFSR_219 :: (IsModule m c) => m (LFSR (Bit 219))
mkLFSR_219 = mkLFSR
mkLFSR_220 :: (IsModule m c) => m (LFSR (Bit 220))
mkLFSR_220 = mkLFSR
mkLFSR_221 :: (IsModule m c) => m (LFSR (Bit 221))
mkLFSR_221 = mkLFSR
mkLFSR_222 :: (IsModule m c) => m (LFSR (Bit 222))
mkLFSR_222 = mkLFSR
mkLFSR_223 :: (IsModule m c) => m (LFSR (Bit 223))
mkLFSR_223 = mkLFSR
mkLFSR_224 :: (IsModule m c) => m (LFSR (Bit 224))
mkLFSR_224 = mkLFSR
mkLFSR_225 :: (IsModule m c) => m (LFSR (Bit 225))
mkLFSR_225 = mkLFSR
mkLFSR_226 :: (IsModule m c) => m (LFSR (Bit 226))
mkLFSR_226 = mkLFSR
mkLFSR_227 :: (IsModule m c) => m (LFSR (Bit 227))
mkLFSR_227 = mkLFSR
mkLFSR_228 :: (IsModule m c) => m (LFSR (Bit 228))
mkLFSR_228 = mkLFSR
mkLFSR_229 :: (IsModule m c) => m (LFSR (Bit 229))
mkLFSR_229 = mkLFSR
mkLFSR_230 :: (IsModule m c) => m (LFSR (Bit 230))
mkLFSR_230 = mkLFSR
mkLFSR_231 :: (IsModule m c) => m (LFSR (Bit 231))
mkLFSR_231 = mkLFSR
mkLFSR_232 :: (IsModule m c) => m (LFSR (Bit 232))
mkLFSR_232 = mkLFSR
mkLFSR_233 :: (IsModule m c) => m (LFSR (Bit 233))
mkLFSR_233 = mkLFSR
mkLFSR_234 :: (IsModule m c) => m (LFSR (Bit 234))
mkLFSR_234 = mkLFSR
mkLFSR_235 :: (IsModule m c) => m (LFSR (Bit 235))
mkLFSR_235 = mkLFSR
mkLFSR_236 :: (IsModule m c) => m (LFSR (Bit 236))
mkLFSR_236 = mkLFSR
mkLFSR_237 :: (IsModule m c) => m (LFSR (Bit 237))
mkLFSR_237 = mkLFSR
mkLFSR_238 :: (IsModule m c) => m (LFSR (Bit 238))
mkLFSR_238 = mkLFSR
mkLFSR_239 :: (IsModule m c) => m (LFSR (Bit 239))
mkLFSR_239 = mkLFSR
mkLFSR_240 :: (IsModule m c) => m (LFSR (Bit 240))
mkLFSR_240 = mkLFSR
mkLFSR_241 :: (IsModule m c) => m (LFSR (Bit 241))
mkLFSR_241 = mkLFSR
mkLFSR_242 :: (IsModule m c) => m (LFSR (Bit 242))
mkLFSR_242 = mkLFSR
mkLFSR_243 :: (IsModule m c) => m (LFSR (Bit 243))
mkLFSR_243 = mkLFSR
mkLFSR_244 :: (IsModule m c) => m (LFSR (Bit 244))
mkLFSR_244 = mkLFSR
mkLFSR_245 :: (IsModule m c) => m (LFSR (Bit 245))
mkLFSR_245 = mkLFSR
mkLFSR_246 :: (IsModule m c) => m (LFSR (Bit 246))
mkLFSR_246 = mkLFSR
mkLFSR_247 :: (IsModule m c) => m (LFSR (Bit 247))
mkLFSR_247 = mkLFSR
mkLFSR_248 :: (IsModule m c) => m (LFSR (Bit 248))
mkLFSR_248 = mkLFSR
mkLFSR_249 :: (IsModule m c) => m (LFSR (Bit 249))
mkLFSR_249 = mkLFSR
mkLFSR_250 :: (IsModule m c) => m (LFSR (Bit 250))
mkLFSR_250 = mkLFSR
mkLFSR_251 :: (IsModule m c) => m (LFSR (Bit 251))
mkLFSR_251 = mkLFSR
mkLFSR_252 :: (IsModule m c) => m (LFSR (Bit 252))
mkLFSR_252 = mkLFSR
mkLFSR_253 :: (IsModule m c) => m (LFSR (Bit 253))
mkLFSR_253 = mkLFSR
mkLFSR_254 :: (IsModule m c) => m (LFSR (Bit 254))
mkLFSR_254 = mkLFSR
mkLFSR_255 :: (IsModule m c) => m (LFSR (Bit 255))
mkLFSR_255 = mkLFSR
mkLFSR_256 :: (IsModule m c) => m (LFSR (Bit 256))
mkLFSR_256 = mkLFSR
mkLFSR_257 :: (IsModule m c) => m (LFSR (Bit 257))
mkLFSR_257 = mkLFSR
mkLFSR_258 :: (IsModule m c) => m (LFSR (Bit 258))
mkLFSR_258 = mkLFSR
mkLFSR_259 :: (IsModule m c) => m (LFSR (Bit 259))
mkLFSR_259 = mkLFSR
mkLFSR_260 :: (IsModule m c) => m (LFSR (Bit 260))
mkLFSR_260 = mkLFSR
mkLFSR_261 :: (IsModule m c) => m (LFSR (Bit 261))
mkLFSR_261 = mkLFSR
mkLFSR_262 :: (IsModule m c) => m (LFSR (Bit 262))
mkLFSR_262 = mkLFSR
mkLFSR_263 :: (IsModule m c) => m (LFSR (Bit 263))
mkLFSR_263 = mkLFSR
mkLFSR_264 :: (IsModule m c) => m (LFSR (Bit 264))
mkLFSR_264 = mkLFSR
mkLFSR_265 :: (IsModule m c) => m (LFSR (Bit 265))
mkLFSR_265 = mkLFSR
mkLFSR_266 :: (IsModule m c) => m (LFSR (Bit 266))
mkLFSR_266 = mkLFSR
mkLFSR_267 :: (IsModule m c) => m (LFSR (Bit 267))
mkLFSR_267 = mkLFSR
mkLFSR_268 :: (IsModule m c) => m (LFSR (Bit 268))
mkLFSR_268 = mkLFSR
mkLFSR_269 :: (IsModule m c) => m (LFSR (Bit 269))
mkLFSR_269 = mkLFSR
mkLFSR_270 :: (IsModule m c) => m (LFSR (Bit 270))
mkLFSR_270 = mkLFSR
mkLFSR_271 :: (IsModule m c) => m (LFSR (Bit 271))
mkLFSR_271 = mkLFSR
mkLFSR_272 :: (IsModule m c) => m (LFSR (Bit 272))
mkLFSR_272 = mkLFSR
mkLFSR_273 :: (IsModule m c) => m (LFSR (Bit 273))
mkLFSR_273 = mkLFSR
mkLFSR_274 :: (IsModule m c) => m (LFSR (Bit 274))
mkLFSR_274 = mkLFSR
mkLFSR_275 :: (IsModule m c) => m (LFSR (Bit 275))
mkLFSR_275 = mkLFSR
mkLFSR_276 :: (IsModule m c) => m (LFSR (Bit 276))
mkLFSR_276 = mkLFSR
mkLFSR_277 :: (IsModule m c) => m (LFSR (Bit 277))
mkLFSR_277 = mkLFSR
mkLFSR_278 :: (IsModule m c) => m (LFSR (Bit 278))
mkLFSR_278 = mkLFSR
mkLFSR_279 :: (IsModule m c) => m (LFSR (Bit 279))
mkLFSR_279 = mkLFSR
mkLFSR_280 :: (IsModule m c) => m (LFSR (Bit 280))
mkLFSR_280 = mkLFSR
mkLFSR_281 :: (IsModule m c) => m (LFSR (Bit 281))
mkLFSR_281 = mkLFSR
mkLFSR_282 :: (IsModule m c) => m (LFSR (Bit 282))
mkLFSR_282 = mkLFSR
mkLFSR_283 :: (IsModule m c) => m (LFSR (Bit 283))
mkLFSR_283 = mkLFSR
mkLFSR_284 :: (IsModule m c) => m (LFSR (Bit 284))
mkLFSR_284 = mkLFSR
mkLFSR_285 :: (IsModule m c) => m (LFSR (Bit 285))
mkLFSR_285 = mkLFSR
mkLFSR_286 :: (IsModule m c) => m (LFSR (Bit 286))
mkLFSR_286 = mkLFSR
mkLFSR_287 :: (IsModule m c) => m (LFSR (Bit 287))
mkLFSR_287 = mkLFSR
mkLFSR_288 :: (IsModule m c) => m (LFSR (Bit 288))
mkLFSR_288 = mkLFSR
mkLFSR_289 :: (IsModule m c) => m (LFSR (Bit 289))
mkLFSR_289 = mkLFSR
mkLFSR_290 :: (IsModule m c) => m (LFSR (Bit 290))
mkLFSR_290 = mkLFSR
mkLFSR_291 :: (IsModule m c) => m (LFSR (Bit 291))
mkLFSR_291 = mkLFSR
mkLFSR_292 :: (IsModule m c) => m (LFSR (Bit 292))
mkLFSR_292 = mkLFSR
mkLFSR_293 :: (IsModule m c) => m (LFSR (Bit 293))
mkLFSR_293 = mkLFSR
mkLFSR_294 :: (IsModule m c) => m (LFSR (Bit 294))
mkLFSR_294 = mkLFSR
mkLFSR_295 :: (IsModule m c) => m (LFSR (Bit 295))
mkLFSR_295 = mkLFSR
mkLFSR_296 :: (IsModule m c) => m (LFSR (Bit 296))
mkLFSR_296 = mkLFSR
mkLFSR_297 :: (IsModule m c) => m (LFSR (Bit 297))
mkLFSR_297 = mkLFSR
mkLFSR_298 :: (IsModule m c) => m (LFSR (Bit 298))
mkLFSR_298 = mkLFSR
mkLFSR_299 :: (IsModule m c) => m (LFSR (Bit 299))
mkLFSR_299 = mkLFSR
mkLFSR_300 :: (IsModule m c) => m (LFSR (Bit 300))
mkLFSR_300 = mkLFSR
mkLFSR_301 :: (IsModule m c) => m (LFSR (Bit 301))
mkLFSR_301 = mkLFSR
mkLFSR_302 :: (IsModule m c) => m (LFSR (Bit 302))
mkLFSR_302 = mkLFSR
mkLFSR_303 :: (IsModule m c) => m (LFSR (Bit 303))
mkLFSR_303 = mkLFSR
mkLFSR_304 :: (IsModule m c) => m (LFSR (Bit 304))
mkLFSR_304 = mkLFSR
mkLFSR_305 :: (IsModule m c) => m (LFSR (Bit 305))
mkLFSR_305 = mkLFSR
mkLFSR_306 :: (IsModule m c) => m (LFSR (Bit 306))
mkLFSR_306 = mkLFSR
mkLFSR_307 :: (IsModule m c) => m (LFSR (Bit 307))
mkLFSR_307 = mkLFSR
mkLFSR_308 :: (IsModule m c) => m (LFSR (Bit 308))
mkLFSR_308 = mkLFSR
mkLFSR_309 :: (IsModule m c) => m (LFSR (Bit 309))
mkLFSR_309 = mkLFSR
mkLFSR_310 :: (IsModule m c) => m (LFSR (Bit 310))
mkLFSR_310 = mkLFSR
mkLFSR_311 :: (IsModule m c) => m (LFSR (Bit 311))
mkLFSR_311 = mkLFSR
mkLFSR_312 :: (IsModule m c) => m (LFSR (Bit 312))
mkLFSR_312 = mkLFSR
mkLFSR_313 :: (IsModule m c) => m (LFSR (Bit 313))
mkLFSR_313 = mkLFSR
mkLFSR_314 :: (IsModule m c) => m (LFSR (Bit 314))
mkLFSR_314 = mkLFSR
mkLFSR_315 :: (IsModule m c) => m (LFSR (Bit 315))
mkLFSR_315 = mkLFSR
mkLFSR_316 :: (IsModule m c) => m (LFSR (Bit 316))
mkLFSR_316 = mkLFSR
mkLFSR_317 :: (IsModule m c) => m (LFSR (Bit 317))
mkLFSR_317 = mkLFSR
mkLFSR_318 :: (IsModule m c) => m (LFSR (Bit 318))
mkLFSR_318 = mkLFSR
mkLFSR_319 :: (IsModule m c) => m (LFSR (Bit 319))
mkLFSR_319 = mkLFSR
mkLFSR_320 :: (IsModule m c) => m (LFSR (Bit 320))
mkLFSR_320 = mkLFSR
mkLFSR_321 :: (IsModule m c) => m (LFSR (Bit 321))
mkLFSR_321 = mkLFSR
mkLFSR_322 :: (IsModule m c) => m (LFSR (Bit 322))
mkLFSR_322 = mkLFSR
mkLFSR_323 :: (IsModule m c) => m (LFSR (Bit 323))
mkLFSR_323 = mkLFSR
mkLFSR_324 :: (IsModule m c) => m (LFSR (Bit 324))
mkLFSR_324 = mkLFSR
mkLFSR_325 :: (IsModule m c) => m (LFSR (Bit 325))
mkLFSR_325 = mkLFSR
mkLFSR_326 :: (IsModule m c) => m (LFSR (Bit 326))
mkLFSR_326 = mkLFSR
mkLFSR_327 :: (IsModule m c) => m (LFSR (Bit 327))
mkLFSR_327 = mkLFSR
mkLFSR_328 :: (IsModule m c) => m (LFSR (Bit 328))
mkLFSR_328 = mkLFSR
mkLFSR_329 :: (IsModule m c) => m (LFSR (Bit 329))
mkLFSR_329 = mkLFSR
mkLFSR_330 :: (IsModule m c) => m (LFSR (Bit 330))
mkLFSR_330 = mkLFSR
mkLFSR_331 :: (IsModule m c) => m (LFSR (Bit 331))
mkLFSR_331 = mkLFSR
mkLFSR_332 :: (IsModule m c) => m (LFSR (Bit 332))
mkLFSR_332 = mkLFSR
mkLFSR_333 :: (IsModule m c) => m (LFSR (Bit 333))
mkLFSR_333 = mkLFSR
mkLFSR_334 :: (IsModule m c) => m (LFSR (Bit 334))
mkLFSR_334 = mkLFSR
mkLFSR_335 :: (IsModule m c) => m (LFSR (Bit 335))
mkLFSR_335 = mkLFSR
mkLFSR_336 :: (IsModule m c) => m (LFSR (Bit 336))
mkLFSR_336 = mkLFSR
mkLFSR_337 :: (IsModule m c) => m (LFSR (Bit 337))
mkLFSR_337 = mkLFSR
mkLFSR_338 :: (IsModule m c) => m (LFSR (Bit 338))
mkLFSR_338 = mkLFSR
mkLFSR_339 :: (IsModule m c) => m (LFSR (Bit 339))
mkLFSR_339 = mkLFSR
mkLFSR_340 :: (IsModule m c) => m (LFSR (Bit 340))
mkLFSR_340 = mkLFSR
mkLFSR_341 :: (IsModule m c) => m (LFSR (Bit 341))
mkLFSR_341 = mkLFSR
mkLFSR_342 :: (IsModule m c) => m (LFSR (Bit 342))
mkLFSR_342 = mkLFSR
mkLFSR_343 :: (IsModule m c) => m (LFSR (Bit 343))
mkLFSR_343 = mkLFSR
mkLFSR_344 :: (IsModule m c) => m (LFSR (Bit 344))
mkLFSR_344 = mkLFSR
mkLFSR_345 :: (IsModule m c) => m (LFSR (Bit 345))
mkLFSR_345 = mkLFSR
mkLFSR_346 :: (IsModule m c) => m (LFSR (Bit 346))
mkLFSR_346 = mkLFSR
mkLFSR_347 :: (IsModule m c) => m (LFSR (Bit 347))
mkLFSR_347 = mkLFSR
mkLFSR_348 :: (IsModule m c) => m (LFSR (Bit 348))
mkLFSR_348 = mkLFSR
mkLFSR_349 :: (IsModule m c) => m (LFSR (Bit 349))
mkLFSR_349 = mkLFSR
mkLFSR_350 :: (IsModule m c) => m (LFSR (Bit 350))
mkLFSR_350 = mkLFSR
mkLFSR_351 :: (IsModule m c) => m (LFSR (Bit 351))
mkLFSR_351 = mkLFSR
mkLFSR_352 :: (IsModule m c) => m (LFSR (Bit 352))
mkLFSR_352 = mkLFSR
mkLFSR_353 :: (IsModule m c) => m (LFSR (Bit 353))
mkLFSR_353 = mkLFSR
mkLFSR_354 :: (IsModule m c) => m (LFSR (Bit 354))
mkLFSR_354 = mkLFSR
mkLFSR_355 :: (IsModule m c) => m (LFSR (Bit 355))
mkLFSR_355 = mkLFSR
mkLFSR_356 :: (IsModule m c) => m (LFSR (Bit 356))
mkLFSR_356 = mkLFSR
mkLFSR_357 :: (IsModule m c) => m (LFSR (Bit 357))
mkLFSR_357 = mkLFSR
mkLFSR_358 :: (IsModule m c) => m (LFSR (Bit 358))
mkLFSR_358 = mkLFSR
mkLFSR_359 :: (IsModule m c) => m (LFSR (Bit 359))
mkLFSR_359 = mkLFSR
mkLFSR_360 :: (IsModule m c) => m (LFSR (Bit 360))
mkLFSR_360 = mkLFSR
mkLFSR_361 :: (IsModule m c) => m (LFSR (Bit 361))
mkLFSR_361 = mkLFSR
mkLFSR_362 :: (IsModule m c) => m (LFSR (Bit 362))
mkLFSR_362 = mkLFSR
mkLFSR_363 :: (IsModule m c) => m (LFSR (Bit 363))
mkLFSR_363 = mkLFSR
mkLFSR_364 :: (IsModule m c) => m (LFSR (Bit 364))
mkLFSR_364 = mkLFSR
mkLFSR_365 :: (IsModule m c) => m (LFSR (Bit 365))
mkLFSR_365 = mkLFSR
mkLFSR_366 :: (IsModule m c) => m (LFSR (Bit 366))
mkLFSR_366 = mkLFSR
mkLFSR_367 :: (IsModule m c) => m (LFSR (Bit 367))
mkLFSR_367 = mkLFSR
mkLFSR_368 :: (IsModule m c) => m (LFSR (Bit 368))
mkLFSR_368 = mkLFSR
mkLFSR_369 :: (IsModule m c) => m (LFSR (Bit 369))
mkLFSR_369 = mkLFSR
mkLFSR_370 :: (IsModule m c) => m (LFSR (Bit 370))
mkLFSR_370 = mkLFSR
mkLFSR_371 :: (IsModule m c) => m (LFSR (Bit 371))
mkLFSR_371 = mkLFSR
mkLFSR_372 :: (IsModule m c) => m (LFSR (Bit 372))
mkLFSR_372 = mkLFSR
mkLFSR_373 :: (IsModule m c) => m (LFSR (Bit 373))
mkLFSR_373 = mkLFSR
mkLFSR_374 :: (IsModule m c) => m (LFSR (Bit 374))
mkLFSR_374 = mkLFSR
mkLFSR_375 :: (IsModule m c) => m (LFSR (Bit 375))
mkLFSR_375 = mkLFSR
mkLFSR_376 :: (IsModule m c) => m (LFSR (Bit 376))
mkLFSR_376 = mkLFSR
mkLFSR_377 :: (IsModule m c) => m (LFSR (Bit 377))
mkLFSR_377 = mkLFSR
mkLFSR_378 :: (IsModule m c) => m (LFSR (Bit 378))
mkLFSR_378 = mkLFSR
mkLFSR_379 :: (IsModule m c) => m (LFSR (Bit 379))
mkLFSR_379 = mkLFSR
mkLFSR_380 :: (IsModule m c) => m (LFSR (Bit 380))
mkLFSR_380 = mkLFSR
mkLFSR_381 :: (IsModule m c) => m (LFSR (Bit 381))
mkLFSR_381 = mkLFSR
mkLFSR_382 :: (IsModule m c) => m (LFSR (Bit 382))
mkLFSR_382 = mkLFSR
mkLFSR_383 :: (IsModule m c) => m (LFSR (Bit 383))
mkLFSR_383 = mkLFSR
mkLFSR_384 :: (IsModule m c) => m (LFSR (Bit 384))
mkLFSR_384 = mkLFSR
mkLFSR_385 :: (IsModule m c) => m (LFSR (Bit 385))
mkLFSR_385 = mkLFSR
mkLFSR_386 :: (IsModule m c) => m (LFSR (Bit 386))
mkLFSR_386 = mkLFSR
mkLFSR_387 :: (IsModule m c) => m (LFSR (Bit 387))
mkLFSR_387 = mkLFSR
mkLFSR_388 :: (IsModule m c) => m (LFSR (Bit 388))
mkLFSR_388 = mkLFSR
mkLFSR_389 :: (IsModule m c) => m (LFSR (Bit 389))
mkLFSR_389 = mkLFSR
mkLFSR_390 :: (IsModule m c) => m (LFSR (Bit 390))
mkLFSR_390 = mkLFSR
mkLFSR_391 :: (IsModule m c) => m (LFSR (Bit 391))
mkLFSR_391 = mkLFSR
mkLFSR_392 :: (IsModule m c) => m (LFSR (Bit 392))
mkLFSR_392 = mkLFSR
mkLFSR_393 :: (IsModule m c) => m (LFSR (Bit 393))
mkLFSR_393 = mkLFSR
mkLFSR_394 :: (IsModule m c) => m (LFSR (Bit 394))
mkLFSR_394 = mkLFSR
mkLFSR_395 :: (IsModule m c) => m (LFSR (Bit 395))
mkLFSR_395 = mkLFSR
mkLFSR_396 :: (IsModule m c) => m (LFSR (Bit 396))
mkLFSR_396 = mkLFSR
mkLFSR_397 :: (IsModule m c) => m (LFSR (Bit 397))
mkLFSR_397 = mkLFSR
mkLFSR_398 :: (IsModule m c) => m (LFSR (Bit 398))
mkLFSR_398 = mkLFSR
mkLFSR_399 :: (IsModule m c) => m (LFSR (Bit 399))
mkLFSR_399 = mkLFSR
mkLFSR_400 :: (IsModule m c) => m (LFSR (Bit 400))
mkLFSR_400 = mkLFSR
mkLFSR_401 :: (IsModule m c) => m (LFSR (Bit 401))
mkLFSR_401 = mkLFSR
mkLFSR_402 :: (IsModule m c) => m (LFSR (Bit 402))
mkLFSR_402 = mkLFSR
mkLFSR_403 :: (IsModule m c) => m (LFSR (Bit 403))
mkLFSR_403 = mkLFSR
mkLFSR_404 :: (IsModule m c) => m (LFSR (Bit 404))
mkLFSR_404 = mkLFSR
mkLFSR_405 :: (IsModule m c) => m (LFSR (Bit 405))
mkLFSR_405 = mkLFSR
mkLFSR_406 :: (IsModule m c) => m (LFSR (Bit 406))
mkLFSR_406 = mkLFSR
mkLFSR_407 :: (IsModule m c) => m (LFSR (Bit 407))
mkLFSR_407 = mkLFSR
mkLFSR_408 :: (IsModule m c) => m (LFSR (Bit 408))
mkLFSR_408 = mkLFSR
mkLFSR_409 :: (IsModule m c) => m (LFSR (Bit 409))
mkLFSR_409 = mkLFSR
mkLFSR_410 :: (IsModule m c) => m (LFSR (Bit 410))
mkLFSR_410 = mkLFSR
mkLFSR_411 :: (IsModule m c) => m (LFSR (Bit 411))
mkLFSR_411 = mkLFSR
mkLFSR_412 :: (IsModule m c) => m (LFSR (Bit 412))
mkLFSR_412 = mkLFSR
mkLFSR_413 :: (IsModule m c) => m (LFSR (Bit 413))
mkLFSR_413 = mkLFSR
mkLFSR_414 :: (IsModule m c) => m (LFSR (Bit 414))
mkLFSR_414 = mkLFSR
mkLFSR_415 :: (IsModule m c) => m (LFSR (Bit 415))
mkLFSR_415 = mkLFSR
mkLFSR_416 :: (IsModule m c) => m (LFSR (Bit 416))
mkLFSR_416 = mkLFSR
mkLFSR_417 :: (IsModule m c) => m (LFSR (Bit 417))
mkLFSR_417 = mkLFSR
mkLFSR_418 :: (IsModule m c) => m (LFSR (Bit 418))
mkLFSR_418 = mkLFSR
mkLFSR_419 :: (IsModule m c) => m (LFSR (Bit 419))
mkLFSR_419 = mkLFSR
mkLFSR_420 :: (IsModule m c) => m (LFSR (Bit 420))
mkLFSR_420 = mkLFSR
mkLFSR_421 :: (IsModule m c) => m (LFSR (Bit 421))
mkLFSR_421 = mkLFSR
mkLFSR_422 :: (IsModule m c) => m (LFSR (Bit 422))
mkLFSR_422 = mkLFSR
mkLFSR_423 :: (IsModule m c) => m (LFSR (Bit 423))
mkLFSR_423 = mkLFSR
mkLFSR_424 :: (IsModule m c) => m (LFSR (Bit 424))
mkLFSR_424 = mkLFSR
mkLFSR_425 :: (IsModule m c) => m (LFSR (Bit 425))
mkLFSR_425 = mkLFSR
mkLFSR_426 :: (IsModule m c) => m (LFSR (Bit 426))
mkLFSR_426 = mkLFSR
mkLFSR_427 :: (IsModule m c) => m (LFSR (Bit 427))
mkLFSR_427 = mkLFSR
mkLFSR_428 :: (IsModule m c) => m (LFSR (Bit 428))
mkLFSR_428 = mkLFSR
mkLFSR_429 :: (IsModule m c) => m (LFSR (Bit 429))
mkLFSR_429 = mkLFSR
mkLFSR_430 :: (IsModule m c) => m (LFSR (Bit 430))
mkLFSR_430 = mkLFSR
mkLFSR_431 :: (IsModule m c) => m (LFSR (Bit 431))
mkLFSR_431 = mkLFSR
mkLFSR_432 :: (IsModule m c) => m (LFSR (Bit 432))
mkLFSR_432 = mkLFSR
mkLFSR_433 :: (IsModule m c) => m (LFSR (Bit 433))
mkLFSR_433 = mkLFSR
mkLFSR_434 :: (IsModule m c) => m (LFSR (Bit 434))
mkLFSR_434 = mkLFSR
mkLFSR_435 :: (IsModule m c) => m (LFSR (Bit 435))
mkLFSR_435 = mkLFSR
mkLFSR_436 :: (IsModule m c) => m (LFSR (Bit 436))
mkLFSR_436 = mkLFSR
mkLFSR_437 :: (IsModule m c) => m (LFSR (Bit 437))
mkLFSR_437 = mkLFSR
mkLFSR_438 :: (IsModule m c) => m (LFSR (Bit 438))
mkLFSR_438 = mkLFSR
mkLFSR_439 :: (IsModule m c) => m (LFSR (Bit 439))
mkLFSR_439 = mkLFSR
mkLFSR_440 :: (IsModule m c) => m (LFSR (Bit 440))
mkLFSR_440 = mkLFSR
mkLFSR_441 :: (IsModule m c) => m (LFSR (Bit 441))
mkLFSR_441 = mkLFSR
mkLFSR_442 :: (IsModule m c) => m (LFSR (Bit 442))
mkLFSR_442 = mkLFSR
mkLFSR_443 :: (IsModule m c) => m (LFSR (Bit 443))
mkLFSR_443 = mkLFSR
mkLFSR_444 :: (IsModule m c) => m (LFSR (Bit 444))
mkLFSR_444 = mkLFSR
mkLFSR_445 :: (IsModule m c) => m (LFSR (Bit 445))
mkLFSR_445 = mkLFSR
mkLFSR_446 :: (IsModule m c) => m (LFSR (Bit 446))
mkLFSR_446 = mkLFSR
mkLFSR_447 :: (IsModule m c) => m (LFSR (Bit 447))
mkLFSR_447 = mkLFSR
mkLFSR_448 :: (IsModule m c) => m (LFSR (Bit 448))
mkLFSR_448 = mkLFSR
mkLFSR_449 :: (IsModule m c) => m (LFSR (Bit 449))
mkLFSR_449 = mkLFSR
mkLFSR_450 :: (IsModule m c) => m (LFSR (Bit 450))
mkLFSR_450 = mkLFSR
mkLFSR_451 :: (IsModule m c) => m (LFSR (Bit 451))
mkLFSR_451 = mkLFSR
mkLFSR_452 :: (IsModule m c) => m (LFSR (Bit 452))
mkLFSR_452 = mkLFSR
mkLFSR_453 :: (IsModule m c) => m (LFSR (Bit 453))
mkLFSR_453 = mkLFSR
mkLFSR_454 :: (IsModule m c) => m (LFSR (Bit 454))
mkLFSR_454 = mkLFSR
mkLFSR_455 :: (IsModule m c) => m (LFSR (Bit 455))
mkLFSR_455 = mkLFSR
mkLFSR_456 :: (IsModule m c) => m (LFSR (Bit 456))
mkLFSR_456 = mkLFSR
mkLFSR_457 :: (IsModule m c) => m (LFSR (Bit 457))
mkLFSR_457 = mkLFSR
mkLFSR_458 :: (IsModule m c) => m (LFSR (Bit 458))
mkLFSR_458 = mkLFSR
mkLFSR_459 :: (IsModule m c) => m (LFSR (Bit 459))
mkLFSR_459 = mkLFSR
mkLFSR_460 :: (IsModule m c) => m (LFSR (Bit 460))
mkLFSR_460 = mkLFSR
mkLFSR_461 :: (IsModule m c) => m (LFSR (Bit 461))
mkLFSR_461 = mkLFSR
mkLFSR_462 :: (IsModule m c) => m (LFSR (Bit 462))
mkLFSR_462 = mkLFSR
mkLFSR_463 :: (IsModule m c) => m (LFSR (Bit 463))
mkLFSR_463 = mkLFSR
mkLFSR_464 :: (IsModule m c) => m (LFSR (Bit 464))
mkLFSR_464 = mkLFSR
mkLFSR_465 :: (IsModule m c) => m (LFSR (Bit 465))
mkLFSR_465 = mkLFSR
mkLFSR_466 :: (IsModule m c) => m (LFSR (Bit 466))
mkLFSR_466 = mkLFSR
mkLFSR_467 :: (IsModule m c) => m (LFSR (Bit 467))
mkLFSR_467 = mkLFSR
mkLFSR_468 :: (IsModule m c) => m (LFSR (Bit 468))
mkLFSR_468 = mkLFSR
mkLFSR_469 :: (IsModule m c) => m (LFSR (Bit 469))
mkLFSR_469 = mkLFSR
mkLFSR_470 :: (IsModule m c) => m (LFSR (Bit 470))
mkLFSR_470 = mkLFSR
mkLFSR_471 :: (IsModule m c) => m (LFSR (Bit 471))
mkLFSR_471 = mkLFSR
mkLFSR_472 :: (IsModule m c) => m (LFSR (Bit 472))
mkLFSR_472 = mkLFSR
mkLFSR_473 :: (IsModule m c) => m (LFSR (Bit 473))
mkLFSR_473 = mkLFSR
mkLFSR_474 :: (IsModule m c) => m (LFSR (Bit 474))
mkLFSR_474 = mkLFSR
mkLFSR_475 :: (IsModule m c) => m (LFSR (Bit 475))
mkLFSR_475 = mkLFSR
mkLFSR_476 :: (IsModule m c) => m (LFSR (Bit 476))
mkLFSR_476 = mkLFSR
mkLFSR_477 :: (IsModule m c) => m (LFSR (Bit 477))
mkLFSR_477 = mkLFSR
mkLFSR_478 :: (IsModule m c) => m (LFSR (Bit 478))
mkLFSR_478 = mkLFSR
mkLFSR_479 :: (IsModule m c) => m (LFSR (Bit 479))
mkLFSR_479 = mkLFSR
mkLFSR_480 :: (IsModule m c) => m (LFSR (Bit 480))
mkLFSR_480 = mkLFSR
mkLFSR_481 :: (IsModule m c) => m (LFSR (Bit 481))
mkLFSR_481 = mkLFSR
mkLFSR_482 :: (IsModule m c) => m (LFSR (Bit 482))
mkLFSR_482 = mkLFSR
mkLFSR_483 :: (IsModule m c) => m (LFSR (Bit 483))
mkLFSR_483 = mkLFSR
mkLFSR_484 :: (IsModule m c) => m (LFSR (Bit 484))
mkLFSR_484 = mkLFSR
mkLFSR_485 :: (IsModule m c) => m (LFSR (Bit 485))
mkLFSR_485 = mkLFSR
mkLFSR_486 :: (IsModule m c) => m (LFSR (Bit 486))
mkLFSR_486 = mkLFSR
mkLFSR_487 :: (IsModule m c) => m (LFSR (Bit 487))
mkLFSR_487 = mkLFSR
mkLFSR_488 :: (IsModule m c) => m (LFSR (Bit 488))
mkLFSR_488 = mkLFSR
mkLFSR_489 :: (IsModule m c) => m (LFSR (Bit 489))
mkLFSR_489 = mkLFSR
mkLFSR_490 :: (IsModule m c) => m (LFSR (Bit 490))
mkLFSR_490 = mkLFSR
mkLFSR_491 :: (IsModule m c) => m (LFSR (Bit 491))
mkLFSR_491 = mkLFSR
mkLFSR_492 :: (IsModule m c) => m (LFSR (Bit 492))
mkLFSR_492 = mkLFSR
mkLFSR_493 :: (IsModule m c) => m (LFSR (Bit 493))
mkLFSR_493 = mkLFSR
mkLFSR_494 :: (IsModule m c) => m (LFSR (Bit 494))
mkLFSR_494 = mkLFSR
mkLFSR_495 :: (IsModule m c) => m (LFSR (Bit 495))
mkLFSR_495 = mkLFSR
mkLFSR_496 :: (IsModule m c) => m (LFSR (Bit 496))
mkLFSR_496 = mkLFSR
mkLFSR_497 :: (IsModule m c) => m (LFSR (Bit 497))
mkLFSR_497 = mkLFSR
mkLFSR_498 :: (IsModule m c) => m (LFSR (Bit 498))
mkLFSR_498 = mkLFSR
mkLFSR_499 :: (IsModule m c) => m (LFSR (Bit 499))
mkLFSR_499 = mkLFSR
mkLFSR_500 :: (IsModule m c) => m (LFSR (Bit 500))
mkLFSR_500 = mkLFSR
mkLFSR_501 :: (IsModule m c) => m (LFSR (Bit 501))
mkLFSR_501 = mkLFSR
mkLFSR_502 :: (IsModule m c) => m (LFSR (Bit 502))
mkLFSR_502 = mkLFSR
mkLFSR_503 :: (IsModule m c) => m (LFSR (Bit 503))
mkLFSR_503 = mkLFSR
mkLFSR_504 :: (IsModule m c) => m (LFSR (Bit 504))
mkLFSR_504 = mkLFSR
mkLFSR_505 :: (IsModule m c) => m (LFSR (Bit 505))
mkLFSR_505 = mkLFSR
mkLFSR_506 :: (IsModule m c) => m (LFSR (Bit 506))
mkLFSR_506 = mkLFSR
mkLFSR_507 :: (IsModule m c) => m (LFSR (Bit 507))
mkLFSR_507 = mkLFSR
mkLFSR_508 :: (IsModule m c) => m (LFSR (Bit 508))
mkLFSR_508 = mkLFSR
mkLFSR_509 :: (IsModule m c) => m (LFSR (Bit 509))
mkLFSR_509 = mkLFSR
mkLFSR_510 :: (IsModule m c) => m (LFSR (Bit 510))
mkLFSR_510 = mkLFSR
mkLFSR_511 :: (IsModule m c) => m (LFSR (Bit 511))
mkLFSR_511 = mkLFSR
mkLFSR_512 :: (IsModule m c) => m (LFSR (Bit 512))
mkLFSR_512 = mkLFSR
mkLFSR_513 :: (IsModule m c) => m (LFSR (Bit 513))
mkLFSR_513 = mkLFSR
mkLFSR_514 :: (IsModule m c) => m (LFSR (Bit 514))
mkLFSR_514 = mkLFSR
mkLFSR_515 :: (IsModule m c) => m (LFSR (Bit 515))
mkLFSR_515 = mkLFSR
mkLFSR_516 :: (IsModule m c) => m (LFSR (Bit 516))
mkLFSR_516 = mkLFSR
mkLFSR_517 :: (IsModule m c) => m (LFSR (Bit 517))
mkLFSR_517 = mkLFSR
mkLFSR_518 :: (IsModule m c) => m (LFSR (Bit 518))
mkLFSR_518 = mkLFSR
mkLFSR_519 :: (IsModule m c) => m (LFSR (Bit 519))
mkLFSR_519 = mkLFSR
mkLFSR_520 :: (IsModule m c) => m (LFSR (Bit 520))
mkLFSR_520 = mkLFSR
mkLFSR_521 :: (IsModule m c) => m (LFSR (Bit 521))
mkLFSR_521 = mkLFSR
mkLFSR_522 :: (IsModule m c) => m (LFSR (Bit 522))
mkLFSR_522 = mkLFSR
mkLFSR_523 :: (IsModule m c) => m (LFSR (Bit 523))
mkLFSR_523 = mkLFSR
mkLFSR_524 :: (IsModule m c) => m (LFSR (Bit 524))
mkLFSR_524 = mkLFSR
mkLFSR_525 :: (IsModule m c) => m (LFSR (Bit 525))
mkLFSR_525 = mkLFSR
mkLFSR_526 :: (IsModule m c) => m (LFSR (Bit 526))
mkLFSR_526 = mkLFSR
mkLFSR_527 :: (IsModule m c) => m (LFSR (Bit 527))
mkLFSR_527 = mkLFSR
mkLFSR_528 :: (IsModule m c) => m (LFSR (Bit 528))
mkLFSR_528 = mkLFSR
mkLFSR_529 :: (IsModule m c) => m (LFSR (Bit 529))
mkLFSR_529 = mkLFSR
mkLFSR_530 :: (IsModule m c) => m (LFSR (Bit 530))
mkLFSR_530 = mkLFSR
mkLFSR_531 :: (IsModule m c) => m (LFSR (Bit 531))
mkLFSR_531 = mkLFSR
mkLFSR_532 :: (IsModule m c) => m (LFSR (Bit 532))
mkLFSR_532 = mkLFSR
mkLFSR_533 :: (IsModule m c) => m (LFSR (Bit 533))
mkLFSR_533 = mkLFSR
mkLFSR_534 :: (IsModule m c) => m (LFSR (Bit 534))
mkLFSR_534 = mkLFSR
mkLFSR_535 :: (IsModule m c) => m (LFSR (Bit 535))
mkLFSR_535 = mkLFSR
mkLFSR_536 :: (IsModule m c) => m (LFSR (Bit 536))
mkLFSR_536 = mkLFSR
mkLFSR_537 :: (IsModule m c) => m (LFSR (Bit 537))
mkLFSR_537 = mkLFSR
mkLFSR_538 :: (IsModule m c) => m (LFSR (Bit 538))
mkLFSR_538 = mkLFSR
mkLFSR_539 :: (IsModule m c) => m (LFSR (Bit 539))
mkLFSR_539 = mkLFSR
mkLFSR_540 :: (IsModule m c) => m (LFSR (Bit 540))
mkLFSR_540 = mkLFSR
mkLFSR_541 :: (IsModule m c) => m (LFSR (Bit 541))
mkLFSR_541 = mkLFSR
mkLFSR_542 :: (IsModule m c) => m (LFSR (Bit 542))
mkLFSR_542 = mkLFSR
mkLFSR_543 :: (IsModule m c) => m (LFSR (Bit 543))
mkLFSR_543 = mkLFSR
mkLFSR_544 :: (IsModule m c) => m (LFSR (Bit 544))
mkLFSR_544 = mkLFSR
mkLFSR_545 :: (IsModule m c) => m (LFSR (Bit 545))
mkLFSR_545 = mkLFSR
mkLFSR_546 :: (IsModule m c) => m (LFSR (Bit 546))
mkLFSR_546 = mkLFSR
mkLFSR_547 :: (IsModule m c) => m (LFSR (Bit 547))
mkLFSR_547 = mkLFSR
mkLFSR_548 :: (IsModule m c) => m (LFSR (Bit 548))
mkLFSR_548 = mkLFSR
mkLFSR_549 :: (IsModule m c) => m (LFSR (Bit 549))
mkLFSR_549 = mkLFSR
mkLFSR_550 :: (IsModule m c) => m (LFSR (Bit 550))
mkLFSR_550 = mkLFSR
mkLFSR_551 :: (IsModule m c) => m (LFSR (Bit 551))
mkLFSR_551 = mkLFSR
mkLFSR_552 :: (IsModule m c) => m (LFSR (Bit 552))
mkLFSR_552 = mkLFSR
mkLFSR_553 :: (IsModule m c) => m (LFSR (Bit 553))
mkLFSR_553 = mkLFSR
mkLFSR_554 :: (IsModule m c) => m (LFSR (Bit 554))
mkLFSR_554 = mkLFSR
mkLFSR_555 :: (IsModule m c) => m (LFSR (Bit 555))
mkLFSR_555 = mkLFSR
mkLFSR_556 :: (IsModule m c) => m (LFSR (Bit 556))
mkLFSR_556 = mkLFSR
mkLFSR_557 :: (IsModule m c) => m (LFSR (Bit 557))
mkLFSR_557 = mkLFSR
mkLFSR_558 :: (IsModule m c) => m (LFSR (Bit 558))
mkLFSR_558 = mkLFSR
mkLFSR_559 :: (IsModule m c) => m (LFSR (Bit 559))
mkLFSR_559 = mkLFSR
mkLFSR_560 :: (IsModule m c) => m (LFSR (Bit 560))
mkLFSR_560 = mkLFSR
mkLFSR_561 :: (IsModule m c) => m (LFSR (Bit 561))
mkLFSR_561 = mkLFSR
mkLFSR_562 :: (IsModule m c) => m (LFSR (Bit 562))
mkLFSR_562 = mkLFSR
mkLFSR_563 :: (IsModule m c) => m (LFSR (Bit 563))
mkLFSR_563 = mkLFSR
mkLFSR_564 :: (IsModule m c) => m (LFSR (Bit 564))
mkLFSR_564 = mkLFSR
mkLFSR_565 :: (IsModule m c) => m (LFSR (Bit 565))
mkLFSR_565 = mkLFSR
mkLFSR_566 :: (IsModule m c) => m (LFSR (Bit 566))
mkLFSR_566 = mkLFSR
mkLFSR_567 :: (IsModule m c) => m (LFSR (Bit 567))
mkLFSR_567 = mkLFSR
mkLFSR_568 :: (IsModule m c) => m (LFSR (Bit 568))
mkLFSR_568 = mkLFSR
mkLFSR_569 :: (IsModule m c) => m (LFSR (Bit 569))
mkLFSR_569 = mkLFSR
mkLFSR_570 :: (IsModule m c) => m (LFSR (Bit 570))
mkLFSR_570 = mkLFSR
mkLFSR_571 :: (IsModule m c) => m (LFSR (Bit 571))
mkLFSR_571 = mkLFSR
mkLFSR_572 :: (IsModule m c) => m (LFSR (Bit 572))
mkLFSR_572 = mkLFSR
mkLFSR_573 :: (IsModule m c) => m (LFSR (Bit 573))
mkLFSR_573 = mkLFSR
mkLFSR_574 :: (IsModule m c) => m (LFSR (Bit 574))
mkLFSR_574 = mkLFSR
mkLFSR_575 :: (IsModule m c) => m (LFSR (Bit 575))
mkLFSR_575 = mkLFSR
mkLFSR_576 :: (IsModule m c) => m (LFSR (Bit 576))
mkLFSR_576 = mkLFSR
mkLFSR_577 :: (IsModule m c) => m (LFSR (Bit 577))
mkLFSR_577 = mkLFSR
mkLFSR_578 :: (IsModule m c) => m (LFSR (Bit 578))
mkLFSR_578 = mkLFSR
mkLFSR_579 :: (IsModule m c) => m (LFSR (Bit 579))
mkLFSR_579 = mkLFSR
mkLFSR_580 :: (IsModule m c) => m (LFSR (Bit 580))
mkLFSR_580 = mkLFSR
mkLFSR_581 :: (IsModule m c) => m (LFSR (Bit 581))
mkLFSR_581 = mkLFSR
mkLFSR_582 :: (IsModule m c) => m (LFSR (Bit 582))
mkLFSR_582 = mkLFSR
mkLFSR_583 :: (IsModule m c) => m (LFSR (Bit 583))
mkLFSR_583 = mkLFSR
mkLFSR_584 :: (IsModule m c) => m (LFSR (Bit 584))
mkLFSR_584 = mkLFSR
mkLFSR_585 :: (IsModule m c) => m (LFSR (Bit 585))
mkLFSR_585 = mkLFSR
mkLFSR_586 :: (IsModule m c) => m (LFSR (Bit 586))
mkLFSR_586 = mkLFSR
mkLFSR_587 :: (IsModule m c) => m (LFSR (Bit 587))
mkLFSR_587 = mkLFSR
mkLFSR_588 :: (IsModule m c) => m (LFSR (Bit 588))
mkLFSR_588 = mkLFSR
mkLFSR_589 :: (IsModule m c) => m (LFSR (Bit 589))
mkLFSR_589 = mkLFSR
mkLFSR_590 :: (IsModule m c) => m (LFSR (Bit 590))
mkLFSR_590 = mkLFSR
mkLFSR_591 :: (IsModule m c) => m (LFSR (Bit 591))
mkLFSR_591 = mkLFSR
mkLFSR_592 :: (IsModule m c) => m (LFSR (Bit 592))
mkLFSR_592 = mkLFSR
mkLFSR_593 :: (IsModule m c) => m (LFSR (Bit 593))
mkLFSR_593 = mkLFSR
mkLFSR_594 :: (IsModule m c) => m (LFSR (Bit 594))
mkLFSR_594 = mkLFSR
mkLFSR_595 :: (IsModule m c) => m (LFSR (Bit 595))
mkLFSR_595 = mkLFSR
mkLFSR_596 :: (IsModule m c) => m (LFSR (Bit 596))
mkLFSR_596 = mkLFSR
mkLFSR_597 :: (IsModule m c) => m (LFSR (Bit 597))
mkLFSR_597 = mkLFSR
mkLFSR_598 :: (IsModule m c) => m (LFSR (Bit 598))
mkLFSR_598 = mkLFSR
mkLFSR_599 :: (IsModule m c) => m (LFSR (Bit 599))
mkLFSR_599 = mkLFSR
mkLFSR_600 :: (IsModule m c) => m (LFSR (Bit 600))
mkLFSR_600 = mkLFSR
mkLFSR_601 :: (IsModule m c) => m (LFSR (Bit 601))
mkLFSR_601 = mkLFSR
mkLFSR_602 :: (IsModule m c) => m (LFSR (Bit 602))
mkLFSR_602 = mkLFSR
mkLFSR_603 :: (IsModule m c) => m (LFSR (Bit 603))
mkLFSR_603 = mkLFSR
mkLFSR_604 :: (IsModule m c) => m (LFSR (Bit 604))
mkLFSR_604 = mkLFSR
mkLFSR_605 :: (IsModule m c) => m (LFSR (Bit 605))
mkLFSR_605 = mkLFSR
mkLFSR_606 :: (IsModule m c) => m (LFSR (Bit 606))
mkLFSR_606 = mkLFSR
mkLFSR_607 :: (IsModule m c) => m (LFSR (Bit 607))
mkLFSR_607 = mkLFSR
mkLFSR_608 :: (IsModule m c) => m (LFSR (Bit 608))
mkLFSR_608 = mkLFSR
mkLFSR_609 :: (IsModule m c) => m (LFSR (Bit 609))
mkLFSR_609 = mkLFSR
mkLFSR_610 :: (IsModule m c) => m (LFSR (Bit 610))
mkLFSR_610 = mkLFSR
mkLFSR_611 :: (IsModule m c) => m (LFSR (Bit 611))
mkLFSR_611 = mkLFSR
mkLFSR_612 :: (IsModule m c) => m (LFSR (Bit 612))
mkLFSR_612 = mkLFSR
mkLFSR_613 :: (IsModule m c) => m (LFSR (Bit 613))
mkLFSR_613 = mkLFSR
mkLFSR_614 :: (IsModule m c) => m (LFSR (Bit 614))
mkLFSR_614 = mkLFSR
mkLFSR_615 :: (IsModule m c) => m (LFSR (Bit 615))
mkLFSR_615 = mkLFSR
mkLFSR_616 :: (IsModule m c) => m (LFSR (Bit 616))
mkLFSR_616 = mkLFSR
mkLFSR_617 :: (IsModule m c) => m (LFSR (Bit 617))
mkLFSR_617 = mkLFSR
mkLFSR_618 :: (IsModule m c) => m (LFSR (Bit 618))
mkLFSR_618 = mkLFSR
mkLFSR_619 :: (IsModule m c) => m (LFSR (Bit 619))
mkLFSR_619 = mkLFSR
mkLFSR_620 :: (IsModule m c) => m (LFSR (Bit 620))
mkLFSR_620 = mkLFSR
mkLFSR_621 :: (IsModule m c) => m (LFSR (Bit 621))
mkLFSR_621 = mkLFSR
mkLFSR_622 :: (IsModule m c) => m (LFSR (Bit 622))
mkLFSR_622 = mkLFSR
mkLFSR_623 :: (IsModule m c) => m (LFSR (Bit 623))
mkLFSR_623 = mkLFSR
mkLFSR_624 :: (IsModule m c) => m (LFSR (Bit 624))
mkLFSR_624 = mkLFSR
mkLFSR_625 :: (IsModule m c) => m (LFSR (Bit 625))
mkLFSR_625 = mkLFSR
mkLFSR_626 :: (IsModule m c) => m (LFSR (Bit 626))
mkLFSR_626 = mkLFSR
mkLFSR_627 :: (IsModule m c) => m (LFSR (Bit 627))
mkLFSR_627 = mkLFSR
mkLFSR_628 :: (IsModule m c) => m (LFSR (Bit 628))
mkLFSR_628 = mkLFSR
mkLFSR_629 :: (IsModule m c) => m (LFSR (Bit 629))
mkLFSR_629 = mkLFSR
mkLFSR_630 :: (IsModule m c) => m (LFSR (Bit 630))
mkLFSR_630 = mkLFSR
mkLFSR_631 :: (IsModule m c) => m (LFSR (Bit 631))
mkLFSR_631 = mkLFSR
mkLFSR_632 :: (IsModule m c) => m (LFSR (Bit 632))
mkLFSR_632 = mkLFSR
mkLFSR_633 :: (IsModule m c) => m (LFSR (Bit 633))
mkLFSR_633 = mkLFSR
mkLFSR_634 :: (IsModule m c) => m (LFSR (Bit 634))
mkLFSR_634 = mkLFSR
mkLFSR_635 :: (IsModule m c) => m (LFSR (Bit 635))
mkLFSR_635 = mkLFSR
mkLFSR_636 :: (IsModule m c) => m (LFSR (Bit 636))
mkLFSR_636 = mkLFSR
mkLFSR_637 :: (IsModule m c) => m (LFSR (Bit 637))
mkLFSR_637 = mkLFSR
mkLFSR_638 :: (IsModule m c) => m (LFSR (Bit 638))
mkLFSR_638 = mkLFSR
mkLFSR_639 :: (IsModule m c) => m (LFSR (Bit 639))
mkLFSR_639 = mkLFSR
mkLFSR_640 :: (IsModule m c) => m (LFSR (Bit 640))
mkLFSR_640 = mkLFSR
mkLFSR_641 :: (IsModule m c) => m (LFSR (Bit 641))
mkLFSR_641 = mkLFSR
mkLFSR_642 :: (IsModule m c) => m (LFSR (Bit 642))
mkLFSR_642 = mkLFSR
mkLFSR_643 :: (IsModule m c) => m (LFSR (Bit 643))
mkLFSR_643 = mkLFSR
mkLFSR_644 :: (IsModule m c) => m (LFSR (Bit 644))
mkLFSR_644 = mkLFSR
mkLFSR_645 :: (IsModule m c) => m (LFSR (Bit 645))
mkLFSR_645 = mkLFSR
mkLFSR_646 :: (IsModule m c) => m (LFSR (Bit 646))
mkLFSR_646 = mkLFSR
mkLFSR_647 :: (IsModule m c) => m (LFSR (Bit 647))
mkLFSR_647 = mkLFSR
mkLFSR_648 :: (IsModule m c) => m (LFSR (Bit 648))
mkLFSR_648 = mkLFSR
mkLFSR_649 :: (IsModule m c) => m (LFSR (Bit 649))
mkLFSR_649 = mkLFSR
mkLFSR_650 :: (IsModule m c) => m (LFSR (Bit 650))
mkLFSR_650 = mkLFSR
mkLFSR_651 :: (IsModule m c) => m (LFSR (Bit 651))
mkLFSR_651 = mkLFSR
mkLFSR_652 :: (IsModule m c) => m (LFSR (Bit 652))
mkLFSR_652 = mkLFSR
mkLFSR_653 :: (IsModule m c) => m (LFSR (Bit 653))
mkLFSR_653 = mkLFSR
mkLFSR_654 :: (IsModule m c) => m (LFSR (Bit 654))
mkLFSR_654 = mkLFSR
mkLFSR_655 :: (IsModule m c) => m (LFSR (Bit 655))
mkLFSR_655 = mkLFSR
mkLFSR_656 :: (IsModule m c) => m (LFSR (Bit 656))
mkLFSR_656 = mkLFSR
mkLFSR_657 :: (IsModule m c) => m (LFSR (Bit 657))
mkLFSR_657 = mkLFSR
mkLFSR_658 :: (IsModule m c) => m (LFSR (Bit 658))
mkLFSR_658 = mkLFSR
mkLFSR_659 :: (IsModule m c) => m (LFSR (Bit 659))
mkLFSR_659 = mkLFSR
mkLFSR_660 :: (IsModule m c) => m (LFSR (Bit 660))
mkLFSR_660 = mkLFSR
mkLFSR_661 :: (IsModule m c) => m (LFSR (Bit 661))
mkLFSR_661 = mkLFSR
mkLFSR_662 :: (IsModule m c) => m (LFSR (Bit 662))
mkLFSR_662 = mkLFSR
mkLFSR_663 :: (IsModule m c) => m (LFSR (Bit 663))
mkLFSR_663 = mkLFSR
mkLFSR_664 :: (IsModule m c) => m (LFSR (Bit 664))
mkLFSR_664 = mkLFSR
mkLFSR_665 :: (IsModule m c) => m (LFSR (Bit 665))
mkLFSR_665 = mkLFSR
mkLFSR_666 :: (IsModule m c) => m (LFSR (Bit 666))
mkLFSR_666 = mkLFSR
mkLFSR_667 :: (IsModule m c) => m (LFSR (Bit 667))
mkLFSR_667 = mkLFSR
mkLFSR_668 :: (IsModule m c) => m (LFSR (Bit 668))
mkLFSR_668 = mkLFSR
mkLFSR_669 :: (IsModule m c) => m (LFSR (Bit 669))
mkLFSR_669 = mkLFSR
mkLFSR_670 :: (IsModule m c) => m (LFSR (Bit 670))
mkLFSR_670 = mkLFSR
mkLFSR_671 :: (IsModule m c) => m (LFSR (Bit 671))
mkLFSR_671 = mkLFSR
mkLFSR_672 :: (IsModule m c) => m (LFSR (Bit 672))
mkLFSR_672 = mkLFSR
mkLFSR_673 :: (IsModule m c) => m (LFSR (Bit 673))
mkLFSR_673 = mkLFSR
mkLFSR_674 :: (IsModule m c) => m (LFSR (Bit 674))
mkLFSR_674 = mkLFSR
mkLFSR_675 :: (IsModule m c) => m (LFSR (Bit 675))
mkLFSR_675 = mkLFSR
mkLFSR_676 :: (IsModule m c) => m (LFSR (Bit 676))
mkLFSR_676 = mkLFSR
mkLFSR_677 :: (IsModule m c) => m (LFSR (Bit 677))
mkLFSR_677 = mkLFSR
mkLFSR_678 :: (IsModule m c) => m (LFSR (Bit 678))
mkLFSR_678 = mkLFSR
mkLFSR_679 :: (IsModule m c) => m (LFSR (Bit 679))
mkLFSR_679 = mkLFSR
mkLFSR_680 :: (IsModule m c) => m (LFSR (Bit 680))
mkLFSR_680 = mkLFSR
mkLFSR_681 :: (IsModule m c) => m (LFSR (Bit 681))
mkLFSR_681 = mkLFSR
mkLFSR_682 :: (IsModule m c) => m (LFSR (Bit 682))
mkLFSR_682 = mkLFSR
mkLFSR_683 :: (IsModule m c) => m (LFSR (Bit 683))
mkLFSR_683 = mkLFSR
mkLFSR_684 :: (IsModule m c) => m (LFSR (Bit 684))
mkLFSR_684 = mkLFSR
mkLFSR_685 :: (IsModule m c) => m (LFSR (Bit 685))
mkLFSR_685 = mkLFSR
mkLFSR_686 :: (IsModule m c) => m (LFSR (Bit 686))
mkLFSR_686 = mkLFSR
mkLFSR_687 :: (IsModule m c) => m (LFSR (Bit 687))
mkLFSR_687 = mkLFSR
mkLFSR_688 :: (IsModule m c) => m (LFSR (Bit 688))
mkLFSR_688 = mkLFSR
mkLFSR_689 :: (IsModule m c) => m (LFSR (Bit 689))
mkLFSR_689 = mkLFSR
mkLFSR_690 :: (IsModule m c) => m (LFSR (Bit 690))
mkLFSR_690 = mkLFSR
mkLFSR_691 :: (IsModule m c) => m (LFSR (Bit 691))
mkLFSR_691 = mkLFSR
mkLFSR_692 :: (IsModule m c) => m (LFSR (Bit 692))
mkLFSR_692 = mkLFSR
mkLFSR_693 :: (IsModule m c) => m (LFSR (Bit 693))
mkLFSR_693 = mkLFSR
mkLFSR_694 :: (IsModule m c) => m (LFSR (Bit 694))
mkLFSR_694 = mkLFSR
mkLFSR_695 :: (IsModule m c) => m (LFSR (Bit 695))
mkLFSR_695 = mkLFSR
mkLFSR_696 :: (IsModule m c) => m (LFSR (Bit 696))
mkLFSR_696 = mkLFSR
mkLFSR_697 :: (IsModule m c) => m (LFSR (Bit 697))
mkLFSR_697 = mkLFSR
mkLFSR_698 :: (IsModule m c) => m (LFSR (Bit 698))
mkLFSR_698 = mkLFSR
mkLFSR_699 :: (IsModule m c) => m (LFSR (Bit 699))
mkLFSR_699 = mkLFSR
mkLFSR_700 :: (IsModule m c) => m (LFSR (Bit 700))
mkLFSR_700 = mkLFSR
mkLFSR_701 :: (IsModule m c) => m (LFSR (Bit 701))
mkLFSR_701 = mkLFSR
mkLFSR_702 :: (IsModule m c) => m (LFSR (Bit 702))
mkLFSR_702 = mkLFSR
mkLFSR_703 :: (IsModule m c) => m (LFSR (Bit 703))
mkLFSR_703 = mkLFSR
mkLFSR_704 :: (IsModule m c) => m (LFSR (Bit 704))
mkLFSR_704 = mkLFSR
mkLFSR_705 :: (IsModule m c) => m (LFSR (Bit 705))
mkLFSR_705 = mkLFSR
mkLFSR_706 :: (IsModule m c) => m (LFSR (Bit 706))
mkLFSR_706 = mkLFSR
mkLFSR_707 :: (IsModule m c) => m (LFSR (Bit 707))
mkLFSR_707 = mkLFSR
mkLFSR_708 :: (IsModule m c) => m (LFSR (Bit 708))
mkLFSR_708 = mkLFSR
mkLFSR_709 :: (IsModule m c) => m (LFSR (Bit 709))
mkLFSR_709 = mkLFSR
mkLFSR_710 :: (IsModule m c) => m (LFSR (Bit 710))
mkLFSR_710 = mkLFSR
mkLFSR_711 :: (IsModule m c) => m (LFSR (Bit 711))
mkLFSR_711 = mkLFSR
mkLFSR_712 :: (IsModule m c) => m (LFSR (Bit 712))
mkLFSR_712 = mkLFSR
mkLFSR_713 :: (IsModule m c) => m (LFSR (Bit 713))
mkLFSR_713 = mkLFSR
mkLFSR_714 :: (IsModule m c) => m (LFSR (Bit 714))
mkLFSR_714 = mkLFSR
mkLFSR_715 :: (IsModule m c) => m (LFSR (Bit 715))
mkLFSR_715 = mkLFSR
mkLFSR_716 :: (IsModule m c) => m (LFSR (Bit 716))
mkLFSR_716 = mkLFSR
mkLFSR_717 :: (IsModule m c) => m (LFSR (Bit 717))
mkLFSR_717 = mkLFSR
mkLFSR_718 :: (IsModule m c) => m (LFSR (Bit 718))
mkLFSR_718 = mkLFSR
mkLFSR_719 :: (IsModule m c) => m (LFSR (Bit 719))
mkLFSR_719 = mkLFSR
mkLFSR_720 :: (IsModule m c) => m (LFSR (Bit 720))
mkLFSR_720 = mkLFSR
mkLFSR_721 :: (IsModule m c) => m (LFSR (Bit 721))
mkLFSR_721 = mkLFSR
mkLFSR_722 :: (IsModule m c) => m (LFSR (Bit 722))
mkLFSR_722 = mkLFSR
mkLFSR_723 :: (IsModule m c) => m (LFSR (Bit 723))
mkLFSR_723 = mkLFSR
mkLFSR_724 :: (IsModule m c) => m (LFSR (Bit 724))
mkLFSR_724 = mkLFSR
mkLFSR_725 :: (IsModule m c) => m (LFSR (Bit 725))
mkLFSR_725 = mkLFSR
mkLFSR_726 :: (IsModule m c) => m (LFSR (Bit 726))
mkLFSR_726 = mkLFSR
mkLFSR_727 :: (IsModule m c) => m (LFSR (Bit 727))
mkLFSR_727 = mkLFSR
mkLFSR_728 :: (IsModule m c) => m (LFSR (Bit 728))
mkLFSR_728 = mkLFSR
mkLFSR_729 :: (IsModule m c) => m (LFSR (Bit 729))
mkLFSR_729 = mkLFSR
mkLFSR_730 :: (IsModule m c) => m (LFSR (Bit 730))
mkLFSR_730 = mkLFSR
mkLFSR_731 :: (IsModule m c) => m (LFSR (Bit 731))
mkLFSR_731 = mkLFSR
mkLFSR_732 :: (IsModule m c) => m (LFSR (Bit 732))
mkLFSR_732 = mkLFSR
mkLFSR_733 :: (IsModule m c) => m (LFSR (Bit 733))
mkLFSR_733 = mkLFSR
mkLFSR_734 :: (IsModule m c) => m (LFSR (Bit 734))
mkLFSR_734 = mkLFSR
mkLFSR_735 :: (IsModule m c) => m (LFSR (Bit 735))
mkLFSR_735 = mkLFSR
mkLFSR_736 :: (IsModule m c) => m (LFSR (Bit 736))
mkLFSR_736 = mkLFSR
mkLFSR_737 :: (IsModule m c) => m (LFSR (Bit 737))
mkLFSR_737 = mkLFSR
mkLFSR_738 :: (IsModule m c) => m (LFSR (Bit 738))
mkLFSR_738 = mkLFSR
mkLFSR_739 :: (IsModule m c) => m (LFSR (Bit 739))
mkLFSR_739 = mkLFSR
mkLFSR_740 :: (IsModule m c) => m (LFSR (Bit 740))
mkLFSR_740 = mkLFSR
mkLFSR_741 :: (IsModule m c) => m (LFSR (Bit 741))
mkLFSR_741 = mkLFSR
mkLFSR_742 :: (IsModule m c) => m (LFSR (Bit 742))
mkLFSR_742 = mkLFSR
mkLFSR_743 :: (IsModule m c) => m (LFSR (Bit 743))
mkLFSR_743 = mkLFSR
mkLFSR_744 :: (IsModule m c) => m (LFSR (Bit 744))
mkLFSR_744 = mkLFSR
mkLFSR_745 :: (IsModule m c) => m (LFSR (Bit 745))
mkLFSR_745 = mkLFSR
mkLFSR_746 :: (IsModule m c) => m (LFSR (Bit 746))
mkLFSR_746 = mkLFSR
mkLFSR_747 :: (IsModule m c) => m (LFSR (Bit 747))
mkLFSR_747 = mkLFSR
mkLFSR_748 :: (IsModule m c) => m (LFSR (Bit 748))
mkLFSR_748 = mkLFSR
mkLFSR_749 :: (IsModule m c) => m (LFSR (Bit 749))
mkLFSR_749 = mkLFSR
mkLFSR_750 :: (IsModule m c) => m (LFSR (Bit 750))
mkLFSR_750 = mkLFSR
mkLFSR_751 :: (IsModule m c) => m (LFSR (Bit 751))
mkLFSR_751 = mkLFSR
mkLFSR_752 :: (IsModule m c) => m (LFSR (Bit 752))
mkLFSR_752 = mkLFSR
mkLFSR_753 :: (IsModule m c) => m (LFSR (Bit 753))
mkLFSR_753 = mkLFSR
mkLFSR_754 :: (IsModule m c) => m (LFSR (Bit 754))
mkLFSR_754 = mkLFSR
mkLFSR_755 :: (IsModule m c) => m (LFSR (Bit 755))
mkLFSR_755 = mkLFSR
mkLFSR_756 :: (IsModule m c) => m (LFSR (Bit 756))
mkLFSR_756 = mkLFSR
mkLFSR_757 :: (IsModule m c) => m (LFSR (Bit 757))
mkLFSR_757 = mkLFSR
mkLFSR_758 :: (IsModule m c) => m (LFSR (Bit 758))
mkLFSR_758 = mkLFSR
mkLFSR_759 :: (IsModule m c) => m (LFSR (Bit 759))
mkLFSR_759 = mkLFSR
mkLFSR_760 :: (IsModule m c) => m (LFSR (Bit 760))
mkLFSR_760 = mkLFSR
mkLFSR_761 :: (IsModule m c) => m (LFSR (Bit 761))
mkLFSR_761 = mkLFSR
mkLFSR_762 :: (IsModule m c) => m (LFSR (Bit 762))
mkLFSR_762 = mkLFSR
mkLFSR_763 :: (IsModule m c) => m (LFSR (Bit 763))
mkLFSR_763 = mkLFSR
mkLFSR_764 :: (IsModule m c) => m (LFSR (Bit 764))
mkLFSR_764 = mkLFSR
mkLFSR_765 :: (IsModule m c) => m (LFSR (Bit 765))
mkLFSR_765 = mkLFSR
mkLFSR_766 :: (IsModule m c) => m (LFSR (Bit 766))
mkLFSR_766 = mkLFSR
mkLFSR_767 :: (IsModule m c) => m (LFSR (Bit 767))
mkLFSR_767 = mkLFSR
mkLFSR_768 :: (IsModule m c) => m (LFSR (Bit 768))
mkLFSR_768 = mkLFSR
mkLFSR_769 :: (IsModule m c) => m (LFSR (Bit 769))
mkLFSR_769 = mkLFSR
mkLFSR_770 :: (IsModule m c) => m (LFSR (Bit 770))
mkLFSR_770 = mkLFSR
mkLFSR_771 :: (IsModule m c) => m (LFSR (Bit 771))
mkLFSR_771 = mkLFSR
mkLFSR_772 :: (IsModule m c) => m (LFSR (Bit 772))
mkLFSR_772 = mkLFSR
mkLFSR_773 :: (IsModule m c) => m (LFSR (Bit 773))
mkLFSR_773 = mkLFSR
mkLFSR_774 :: (IsModule m c) => m (LFSR (Bit 774))
mkLFSR_774 = mkLFSR
mkLFSR_775 :: (IsModule m c) => m (LFSR (Bit 775))
mkLFSR_775 = mkLFSR
mkLFSR_776 :: (IsModule m c) => m (LFSR (Bit 776))
mkLFSR_776 = mkLFSR
mkLFSR_777 :: (IsModule m c) => m (LFSR (Bit 777))
mkLFSR_777 = mkLFSR
mkLFSR_778 :: (IsModule m c) => m (LFSR (Bit 778))
mkLFSR_778 = mkLFSR
mkLFSR_779 :: (IsModule m c) => m (LFSR (Bit 779))
mkLFSR_779 = mkLFSR
mkLFSR_780 :: (IsModule m c) => m (LFSR (Bit 780))
mkLFSR_780 = mkLFSR
mkLFSR_781 :: (IsModule m c) => m (LFSR (Bit 781))
mkLFSR_781 = mkLFSR
mkLFSR_782 :: (IsModule m c) => m (LFSR (Bit 782))
mkLFSR_782 = mkLFSR
mkLFSR_783 :: (IsModule m c) => m (LFSR (Bit 783))
mkLFSR_783 = mkLFSR
mkLFSR_784 :: (IsModule m c) => m (LFSR (Bit 784))
mkLFSR_784 = mkLFSR
mkLFSR_785 :: (IsModule m c) => m (LFSR (Bit 785))
mkLFSR_785 = mkLFSR
mkLFSR_786 :: (IsModule m c) => m (LFSR (Bit 786))
mkLFSR_786 = mkLFSR
mkLFSR_787 :: (IsModule m c) => m (LFSR (Bit 787))
mkLFSR_787 = mkLFSR
mkLFSR_788 :: (IsModule m c) => m (LFSR (Bit 788))
mkLFSR_788 = mkLFSR
mkLFSR_789 :: (IsModule m c) => m (LFSR (Bit 789))
mkLFSR_789 = mkLFSR
mkLFSR_790 :: (IsModule m c) => m (LFSR (Bit 790))
mkLFSR_790 = mkLFSR
mkLFSR_791 :: (IsModule m c) => m (LFSR (Bit 791))
mkLFSR_791 = mkLFSR
mkLFSR_792 :: (IsModule m c) => m (LFSR (Bit 792))
mkLFSR_792 = mkLFSR
mkLFSR_793 :: (IsModule m c) => m (LFSR (Bit 793))
mkLFSR_793 = mkLFSR
mkLFSR_794 :: (IsModule m c) => m (LFSR (Bit 794))
mkLFSR_794 = mkLFSR
mkLFSR_795 :: (IsModule m c) => m (LFSR (Bit 795))
mkLFSR_795 = mkLFSR
mkLFSR_796 :: (IsModule m c) => m (LFSR (Bit 796))
mkLFSR_796 = mkLFSR
mkLFSR_797 :: (IsModule m c) => m (LFSR (Bit 797))
mkLFSR_797 = mkLFSR
mkLFSR_798 :: (IsModule m c) => m (LFSR (Bit 798))
mkLFSR_798 = mkLFSR
mkLFSR_799 :: (IsModule m c) => m (LFSR (Bit 799))
mkLFSR_799 = mkLFSR
mkLFSR_800 :: (IsModule m c) => m (LFSR (Bit 800))
mkLFSR_800 = mkLFSR
mkLFSR_801 :: (IsModule m c) => m (LFSR (Bit 801))
mkLFSR_801 = mkLFSR
mkLFSR_802 :: (IsModule m c) => m (LFSR (Bit 802))
mkLFSR_802 = mkLFSR
mkLFSR_803 :: (IsModule m c) => m (LFSR (Bit 803))
mkLFSR_803 = mkLFSR
mkLFSR_804 :: (IsModule m c) => m (LFSR (Bit 804))
mkLFSR_804 = mkLFSR
mkLFSR_805 :: (IsModule m c) => m (LFSR (Bit 805))
mkLFSR_805 = mkLFSR
mkLFSR_806 :: (IsModule m c) => m (LFSR (Bit 806))
mkLFSR_806 = mkLFSR
mkLFSR_807 :: (IsModule m c) => m (LFSR (Bit 807))
mkLFSR_807 = mkLFSR
mkLFSR_808 :: (IsModule m c) => m (LFSR (Bit 808))
mkLFSR_808 = mkLFSR
mkLFSR_809 :: (IsModule m c) => m (LFSR (Bit 809))
mkLFSR_809 = mkLFSR
mkLFSR_810 :: (IsModule m c) => m (LFSR (Bit 810))
mkLFSR_810 = mkLFSR
mkLFSR_811 :: (IsModule m c) => m (LFSR (Bit 811))
mkLFSR_811 = mkLFSR
mkLFSR_812 :: (IsModule m c) => m (LFSR (Bit 812))
mkLFSR_812 = mkLFSR
mkLFSR_813 :: (IsModule m c) => m (LFSR (Bit 813))
mkLFSR_813 = mkLFSR
mkLFSR_814 :: (IsModule m c) => m (LFSR (Bit 814))
mkLFSR_814 = mkLFSR
mkLFSR_815 :: (IsModule m c) => m (LFSR (Bit 815))
mkLFSR_815 = mkLFSR
mkLFSR_816 :: (IsModule m c) => m (LFSR (Bit 816))
mkLFSR_816 = mkLFSR
mkLFSR_817 :: (IsModule m c) => m (LFSR (Bit 817))
mkLFSR_817 = mkLFSR
mkLFSR_818 :: (IsModule m c) => m (LFSR (Bit 818))
mkLFSR_818 = mkLFSR
mkLFSR_819 :: (IsModule m c) => m (LFSR (Bit 819))
mkLFSR_819 = mkLFSR
mkLFSR_820 :: (IsModule m c) => m (LFSR (Bit 820))
mkLFSR_820 = mkLFSR
mkLFSR_821 :: (IsModule m c) => m (LFSR (Bit 821))
mkLFSR_821 = mkLFSR
mkLFSR_822 :: (IsModule m c) => m (LFSR (Bit 822))
mkLFSR_822 = mkLFSR
mkLFSR_823 :: (IsModule m c) => m (LFSR (Bit 823))
mkLFSR_823 = mkLFSR
mkLFSR_824 :: (IsModule m c) => m (LFSR (Bit 824))
mkLFSR_824 = mkLFSR
mkLFSR_825 :: (IsModule m c) => m (LFSR (Bit 825))
mkLFSR_825 = mkLFSR
mkLFSR_826 :: (IsModule m c) => m (LFSR (Bit 826))
mkLFSR_826 = mkLFSR
mkLFSR_827 :: (IsModule m c) => m (LFSR (Bit 827))
mkLFSR_827 = mkLFSR
mkLFSR_828 :: (IsModule m c) => m (LFSR (Bit 828))
mkLFSR_828 = mkLFSR
mkLFSR_829 :: (IsModule m c) => m (LFSR (Bit 829))
mkLFSR_829 = mkLFSR
mkLFSR_830 :: (IsModule m c) => m (LFSR (Bit 830))
mkLFSR_830 = mkLFSR
mkLFSR_831 :: (IsModule m c) => m (LFSR (Bit 831))
mkLFSR_831 = mkLFSR
mkLFSR_832 :: (IsModule m c) => m (LFSR (Bit 832))
mkLFSR_832 = mkLFSR
mkLFSR_833 :: (IsModule m c) => m (LFSR (Bit 833))
mkLFSR_833 = mkLFSR
mkLFSR_834 :: (IsModule m c) => m (LFSR (Bit 834))
mkLFSR_834 = mkLFSR
mkLFSR_835 :: (IsModule m c) => m (LFSR (Bit 835))
mkLFSR_835 = mkLFSR
mkLFSR_836 :: (IsModule m c) => m (LFSR (Bit 836))
mkLFSR_836 = mkLFSR
mkLFSR_837 :: (IsModule m c) => m (LFSR (Bit 837))
mkLFSR_837 = mkLFSR
mkLFSR_838 :: (IsModule m c) => m (LFSR (Bit 838))
mkLFSR_838 = mkLFSR
mkLFSR_839 :: (IsModule m c) => m (LFSR (Bit 839))
mkLFSR_839 = mkLFSR
mkLFSR_840 :: (IsModule m c) => m (LFSR (Bit 840))
mkLFSR_840 = mkLFSR
mkLFSR_841 :: (IsModule m c) => m (LFSR (Bit 841))
mkLFSR_841 = mkLFSR
mkLFSR_842 :: (IsModule m c) => m (LFSR (Bit 842))
mkLFSR_842 = mkLFSR
mkLFSR_843 :: (IsModule m c) => m (LFSR (Bit 843))
mkLFSR_843 = mkLFSR
mkLFSR_844 :: (IsModule m c) => m (LFSR (Bit 844))
mkLFSR_844 = mkLFSR
mkLFSR_845 :: (IsModule m c) => m (LFSR (Bit 845))
mkLFSR_845 = mkLFSR
mkLFSR_846 :: (IsModule m c) => m (LFSR (Bit 846))
mkLFSR_846 = mkLFSR
mkLFSR_847 :: (IsModule m c) => m (LFSR (Bit 847))
mkLFSR_847 = mkLFSR
mkLFSR_848 :: (IsModule m c) => m (LFSR (Bit 848))
mkLFSR_848 = mkLFSR
mkLFSR_849 :: (IsModule m c) => m (LFSR (Bit 849))
mkLFSR_849 = mkLFSR
mkLFSR_850 :: (IsModule m c) => m (LFSR (Bit 850))
mkLFSR_850 = mkLFSR
mkLFSR_851 :: (IsModule m c) => m (LFSR (Bit 851))
mkLFSR_851 = mkLFSR
mkLFSR_852 :: (IsModule m c) => m (LFSR (Bit 852))
mkLFSR_852 = mkLFSR
mkLFSR_853 :: (IsModule m c) => m (LFSR (Bit 853))
mkLFSR_853 = mkLFSR
mkLFSR_854 :: (IsModule m c) => m (LFSR (Bit 854))
mkLFSR_854 = mkLFSR
mkLFSR_855 :: (IsModule m c) => m (LFSR (Bit 855))
mkLFSR_855 = mkLFSR
mkLFSR_856 :: (IsModule m c) => m (LFSR (Bit 856))
mkLFSR_856 = mkLFSR
mkLFSR_857 :: (IsModule m c) => m (LFSR (Bit 857))
mkLFSR_857 = mkLFSR
mkLFSR_858 :: (IsModule m c) => m (LFSR (Bit 858))
mkLFSR_858 = mkLFSR
mkLFSR_859 :: (IsModule m c) => m (LFSR (Bit 859))
mkLFSR_859 = mkLFSR
mkLFSR_860 :: (IsModule m c) => m (LFSR (Bit 860))
mkLFSR_860 = mkLFSR
mkLFSR_861 :: (IsModule m c) => m (LFSR (Bit 861))
mkLFSR_861 = mkLFSR
mkLFSR_862 :: (IsModule m c) => m (LFSR (Bit 862))
mkLFSR_862 = mkLFSR
mkLFSR_863 :: (IsModule m c) => m (LFSR (Bit 863))
mkLFSR_863 = mkLFSR
mkLFSR_864 :: (IsModule m c) => m (LFSR (Bit 864))
mkLFSR_864 = mkLFSR
mkLFSR_865 :: (IsModule m c) => m (LFSR (Bit 865))
mkLFSR_865 = mkLFSR
mkLFSR_866 :: (IsModule m c) => m (LFSR (Bit 866))
mkLFSR_866 = mkLFSR
mkLFSR_867 :: (IsModule m c) => m (LFSR (Bit 867))
mkLFSR_867 = mkLFSR
mkLFSR_868 :: (IsModule m c) => m (LFSR (Bit 868))
mkLFSR_868 = mkLFSR
mkLFSR_869 :: (IsModule m c) => m (LFSR (Bit 869))
mkLFSR_869 = mkLFSR
mkLFSR_870 :: (IsModule m c) => m (LFSR (Bit 870))
mkLFSR_870 = mkLFSR
mkLFSR_871 :: (IsModule m c) => m (LFSR (Bit 871))
mkLFSR_871 = mkLFSR
mkLFSR_872 :: (IsModule m c) => m (LFSR (Bit 872))
mkLFSR_872 = mkLFSR
mkLFSR_873 :: (IsModule m c) => m (LFSR (Bit 873))
mkLFSR_873 = mkLFSR
mkLFSR_874 :: (IsModule m c) => m (LFSR (Bit 874))
mkLFSR_874 = mkLFSR
mkLFSR_875 :: (IsModule m c) => m (LFSR (Bit 875))
mkLFSR_875 = mkLFSR
mkLFSR_876 :: (IsModule m c) => m (LFSR (Bit 876))
mkLFSR_876 = mkLFSR
mkLFSR_877 :: (IsModule m c) => m (LFSR (Bit 877))
mkLFSR_877 = mkLFSR
mkLFSR_878 :: (IsModule m c) => m (LFSR (Bit 878))
mkLFSR_878 = mkLFSR
mkLFSR_879 :: (IsModule m c) => m (LFSR (Bit 879))
mkLFSR_879 = mkLFSR
mkLFSR_880 :: (IsModule m c) => m (LFSR (Bit 880))
mkLFSR_880 = mkLFSR
mkLFSR_881 :: (IsModule m c) => m (LFSR (Bit 881))
mkLFSR_881 = mkLFSR
mkLFSR_882 :: (IsModule m c) => m (LFSR (Bit 882))
mkLFSR_882 = mkLFSR
mkLFSR_883 :: (IsModule m c) => m (LFSR (Bit 883))
mkLFSR_883 = mkLFSR
mkLFSR_884 :: (IsModule m c) => m (LFSR (Bit 884))
mkLFSR_884 = mkLFSR
mkLFSR_885 :: (IsModule m c) => m (LFSR (Bit 885))
mkLFSR_885 = mkLFSR
mkLFSR_886 :: (IsModule m c) => m (LFSR (Bit 886))
mkLFSR_886 = mkLFSR
mkLFSR_887 :: (IsModule m c) => m (LFSR (Bit 887))
mkLFSR_887 = mkLFSR
mkLFSR_888 :: (IsModule m c) => m (LFSR (Bit 888))
mkLFSR_888 = mkLFSR
mkLFSR_889 :: (IsModule m c) => m (LFSR (Bit 889))
mkLFSR_889 = mkLFSR
mkLFSR_890 :: (IsModule m c) => m (LFSR (Bit 890))
mkLFSR_890 = mkLFSR
mkLFSR_891 :: (IsModule m c) => m (LFSR (Bit 891))
mkLFSR_891 = mkLFSR
mkLFSR_892 :: (IsModule m c) => m (LFSR (Bit 892))
mkLFSR_892 = mkLFSR
mkLFSR_893 :: (IsModule m c) => m (LFSR (Bit 893))
mkLFSR_893 = mkLFSR
mkLFSR_894 :: (IsModule m c) => m (LFSR (Bit 894))
mkLFSR_894 = mkLFSR
mkLFSR_895 :: (IsModule m c) => m (LFSR (Bit 895))
mkLFSR_895 = mkLFSR
mkLFSR_896 :: (IsModule m c) => m (LFSR (Bit 896))
mkLFSR_896 = mkLFSR
mkLFSR_897 :: (IsModule m c) => m (LFSR (Bit 897))
mkLFSR_897 = mkLFSR
mkLFSR_898 :: (IsModule m c) => m (LFSR (Bit 898))
mkLFSR_898 = mkLFSR
mkLFSR_899 :: (IsModule m c) => m (LFSR (Bit 899))
mkLFSR_899 = mkLFSR
mkLFSR_900 :: (IsModule m c) => m (LFSR (Bit 900))
mkLFSR_900 = mkLFSR
mkLFSR_901 :: (IsModule m c) => m (LFSR (Bit 901))
mkLFSR_901 = mkLFSR
mkLFSR_902 :: (IsModule m c) => m (LFSR (Bit 902))
mkLFSR_902 = mkLFSR
mkLFSR_903 :: (IsModule m c) => m (LFSR (Bit 903))
mkLFSR_903 = mkLFSR
mkLFSR_904 :: (IsModule m c) => m (LFSR (Bit 904))
mkLFSR_904 = mkLFSR
mkLFSR_905 :: (IsModule m c) => m (LFSR (Bit 905))
mkLFSR_905 = mkLFSR
mkLFSR_906 :: (IsModule m c) => m (LFSR (Bit 906))
mkLFSR_906 = mkLFSR
mkLFSR_907 :: (IsModule m c) => m (LFSR (Bit 907))
mkLFSR_907 = mkLFSR
mkLFSR_908 :: (IsModule m c) => m (LFSR (Bit 908))
mkLFSR_908 = mkLFSR
mkLFSR_909 :: (IsModule m c) => m (LFSR (Bit 909))
mkLFSR_909 = mkLFSR
mkLFSR_910 :: (IsModule m c) => m (LFSR (Bit 910))
mkLFSR_910 = mkLFSR
mkLFSR_911 :: (IsModule m c) => m (LFSR (Bit 911))
mkLFSR_911 = mkLFSR
mkLFSR_912 :: (IsModule m c) => m (LFSR (Bit 912))
mkLFSR_912 = mkLFSR
mkLFSR_913 :: (IsModule m c) => m (LFSR (Bit 913))
mkLFSR_913 = mkLFSR
mkLFSR_914 :: (IsModule m c) => m (LFSR (Bit 914))
mkLFSR_914 = mkLFSR
mkLFSR_915 :: (IsModule m c) => m (LFSR (Bit 915))
mkLFSR_915 = mkLFSR
mkLFSR_916 :: (IsModule m c) => m (LFSR (Bit 916))
mkLFSR_916 = mkLFSR
mkLFSR_917 :: (IsModule m c) => m (LFSR (Bit 917))
mkLFSR_917 = mkLFSR
mkLFSR_918 :: (IsModule m c) => m (LFSR (Bit 918))
mkLFSR_918 = mkLFSR
mkLFSR_919 :: (IsModule m c) => m (LFSR (Bit 919))
mkLFSR_919 = mkLFSR
mkLFSR_920 :: (IsModule m c) => m (LFSR (Bit 920))
mkLFSR_920 = mkLFSR
mkLFSR_921 :: (IsModule m c) => m (LFSR (Bit 921))
mkLFSR_921 = mkLFSR
mkLFSR_922 :: (IsModule m c) => m (LFSR (Bit 922))
mkLFSR_922 = mkLFSR
mkLFSR_923 :: (IsModule m c) => m (LFSR (Bit 923))
mkLFSR_923 = mkLFSR
mkLFSR_924 :: (IsModule m c) => m (LFSR (Bit 924))
mkLFSR_924 = mkLFSR
mkLFSR_925 :: (IsModule m c) => m (LFSR (Bit 925))
mkLFSR_925 = mkLFSR
mkLFSR_926 :: (IsModule m c) => m (LFSR (Bit 926))
mkLFSR_926 = mkLFSR
mkLFSR_927 :: (IsModule m c) => m (LFSR (Bit 927))
mkLFSR_927 = mkLFSR
mkLFSR_928 :: (IsModule m c) => m (LFSR (Bit 928))
mkLFSR_928 = mkLFSR

-- This typeclass lets you generate large random values by combining multiple
-- smaller LFSRs together.

mkRandom :: (IsModule m c, Bits t n, Random n) => m t
mkRandom = mkRandomN 0

class Random n where
  mkRandomN :: (IsModule m c, Bits t n) => Integer -> m t

-- The a and b values of the leaf-nodes of the recursion will "probably not be
-- the same" as each other which is a nice-to-have (but not required) property.
-- This generic instance only kicks in when n is greater then the longest
-- polynomial we have defined, so n//3 will still be "pretty darn big".
instance (Div n 3 d, Add d 7 a,  -- a = n//3 + 7
          Add a b n,             -- b = n - a  (Whatever is left)
          Random a, Random b) => Random n where
  mkRandomN i = module
    a :: Bit a <- mkRandomN (i + 5)
    b :: Bit b <- mkRandomN (i + 3)
    return $ unpack $ a ++ b

-- The explicit instances for the "leaf" LFSRs.
instance Random 2 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 3 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 4 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 5 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 6 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 7 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 8 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 9 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 10 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 11 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 12 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 13 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 14 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 15 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 16 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 17 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 18 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 19 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 20 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 21 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 22 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 23 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 24 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 25 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 26 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 27 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 28 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 29 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 30 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 31 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 32 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 33 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 34 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 35 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 36 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 37 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 38 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 39 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 40 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 41 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 42 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 43 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 44 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 45 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 46 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 47 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 48 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 49 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 50 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 51 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 52 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 53 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 54 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 55 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 56 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 57 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 58 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 59 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 60 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 61 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 62 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 63 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 64 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 65 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 66 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 67 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 68 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 69 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 70 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 71 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 72 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 73 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 74 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 75 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 76 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 77 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 78 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 79 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 80 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 81 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 82 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 83 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 84 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 85 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 86 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 87 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 88 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 89 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 90 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 91 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 92 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 93 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 94 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 95 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 96 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 97 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 98 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 99 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 100 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 101 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 102 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 103 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 104 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 105 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 106 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 107 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 108 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 109 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 110 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 111 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 112 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 113 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 114 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 115 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 116 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 117 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 118 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 119 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 120 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 121 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 122 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 123 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 124 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 125 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 126 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 127 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 128 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 129 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 130 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 131 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 132 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 133 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 134 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 135 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 136 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 137 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 138 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 139 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 140 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 141 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 142 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 143 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 144 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 145 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 146 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 147 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 148 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 149 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 150 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 151 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 152 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 153 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 154 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 155 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 156 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 157 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 158 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 159 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 160 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 161 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 162 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 163 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 164 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 165 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 166 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 167 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 168 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 169 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 170 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 171 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 172 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 173 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 174 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 175 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 176 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 177 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 178 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 179 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 180 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 181 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 182 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 183 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 184 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 185 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 186 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 187 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 188 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 189 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 190 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 191 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 192 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 193 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 194 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 195 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 196 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 197 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 198 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 199 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 200 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 201 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 202 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 203 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 204 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 205 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 206 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 207 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 208 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 209 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 210 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 211 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 212 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 213 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 214 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 215 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 216 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 217 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 218 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 219 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 220 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 221 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 222 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 223 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 224 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 225 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 226 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 227 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 228 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 229 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 230 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 231 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 232 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 233 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 234 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 235 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 236 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 237 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 238 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 239 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 240 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 241 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 242 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 243 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 244 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 245 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 246 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 247 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 248 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 249 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 250 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 251 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 252 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 253 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 254 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 255 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 256 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 257 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 258 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 259 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 260 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 261 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 262 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 263 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 264 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 265 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 266 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 267 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 268 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 269 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 270 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 271 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 272 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 273 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 274 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 275 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 276 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 277 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 278 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 279 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 280 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 281 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 282 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 283 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 284 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 285 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 286 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 287 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 288 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 289 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 290 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 291 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 292 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 293 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 294 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 295 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 296 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 297 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 298 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 299 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 300 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 301 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 302 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 303 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 304 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 305 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 306 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 307 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 308 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 309 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 310 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 311 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 312 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 313 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 314 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 315 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 316 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 317 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 318 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 319 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 320 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 321 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 322 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 323 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 324 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 325 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 326 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 327 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 328 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 329 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 330 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 331 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 332 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 333 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 334 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 335 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 336 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 337 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 338 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 339 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 340 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 341 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 342 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 343 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 344 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 345 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 346 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 347 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 348 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 349 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 350 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 351 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 352 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 353 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 354 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 355 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 356 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 357 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 358 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 359 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 360 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 361 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 362 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 363 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 364 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 365 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 366 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 367 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 368 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 369 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 370 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 371 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 372 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 373 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 374 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 375 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 376 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 377 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 378 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 379 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 380 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 381 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 382 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 383 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 384 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 385 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 386 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 387 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 388 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 389 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 390 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 391 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 392 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 393 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 394 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 395 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 396 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 397 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 398 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 399 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 400 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 401 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 402 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 403 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 404 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 405 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 406 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 407 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 408 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 409 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 410 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 411 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 412 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 413 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 414 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 415 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 416 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 417 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 418 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 419 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 420 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 421 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 422 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 423 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 424 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 425 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 426 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 427 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 428 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 429 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 430 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 431 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 432 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 433 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 434 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 435 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 436 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 437 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 438 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 439 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 440 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 441 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 442 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 443 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 444 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 445 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 446 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 447 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 448 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 449 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 450 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 451 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 452 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 453 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 454 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 455 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 456 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 457 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 458 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 459 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 460 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 461 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 462 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 463 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 464 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 465 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 466 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 467 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 468 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 469 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 470 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 471 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 472 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 473 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 474 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 475 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 476 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 477 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 478 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 479 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 480 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 481 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 482 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 483 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 484 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 485 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 486 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 487 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 488 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 489 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 490 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 491 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 492 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 493 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 494 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 495 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 496 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 497 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 498 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 499 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 500 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 501 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 502 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 503 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 504 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 505 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 506 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 507 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 508 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 509 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 510 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 511 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 512 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 513 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 514 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 515 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 516 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 517 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 518 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 519 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 520 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 521 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 522 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 523 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 524 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 525 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 526 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 527 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 528 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 529 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 530 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 531 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 532 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 533 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 534 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 535 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 536 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 537 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 538 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 539 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 540 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 541 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 542 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 543 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 544 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 545 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 546 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 547 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 548 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 549 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 550 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 551 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 552 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 553 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 554 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 555 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 556 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 557 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 558 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 559 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 560 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 561 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 562 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 563 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 564 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 565 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 566 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 567 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 568 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 569 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 570 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 571 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 572 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 573 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 574 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 575 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 576 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 577 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 578 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 579 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 580 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 581 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 582 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 583 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 584 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 585 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 586 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 587 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 588 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 589 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 590 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 591 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 592 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 593 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 594 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 595 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 596 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 597 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 598 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 599 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 600 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 601 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 602 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 603 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 604 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 605 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 606 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 607 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 608 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 609 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 610 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 611 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 612 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 613 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 614 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 615 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 616 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 617 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 618 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 619 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 620 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 621 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 622 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 623 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 624 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 625 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 626 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 627 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 628 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 629 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 630 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 631 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 632 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 633 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 634 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 635 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 636 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 637 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 638 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 639 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 640 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 641 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 642 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 643 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 644 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 645 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 646 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 647 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 648 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 649 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 650 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 651 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 652 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 653 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 654 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 655 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 656 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 657 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 658 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 659 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 660 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 661 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 662 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 663 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 664 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 665 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 666 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 667 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 668 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 669 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 670 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 671 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 672 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 673 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 674 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 675 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 676 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 677 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 678 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 679 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 680 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 681 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 682 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 683 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 684 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 685 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 686 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 687 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 688 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 689 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 690 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 691 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 692 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 693 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 694 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 695 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 696 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 697 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 698 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 699 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 700 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 701 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 702 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 703 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 704 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 705 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 706 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 707 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 708 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 709 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 710 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 711 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 712 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 713 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 714 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 715 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 716 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 717 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 718 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 719 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 720 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 721 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 722 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 723 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 724 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 725 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 726 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 727 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 728 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 729 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 730 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 731 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 732 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 733 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 734 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 735 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 736 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 737 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 738 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 739 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 740 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 741 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 742 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 743 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 744 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 745 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 746 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 747 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 748 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 749 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 750 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 751 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 752 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 753 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 754 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 755 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 756 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 757 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 758 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 759 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 760 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 761 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 762 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 763 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 764 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 765 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 766 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 767 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 768 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 769 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 770 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 771 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 772 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 773 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 774 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 775 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 776 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 777 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 778 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 779 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 780 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 781 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 782 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 783 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 784 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 785 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 786 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 787 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 788 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 789 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 790 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 791 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 792 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 793 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 794 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 795 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 796 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 797 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 798 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 799 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 800 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 801 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 802 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 803 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 804 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 805 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 806 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 807 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 808 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 809 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 810 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 811 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 812 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 813 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 814 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 815 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 816 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 817 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 818 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 819 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 820 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 821 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 822 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 823 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 824 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 825 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 826 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 827 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 828 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 829 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 830 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 831 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 832 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 833 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 834 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 835 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 836 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 837 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 838 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 839 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 840 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 841 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 842 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 843 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 844 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 845 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 846 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 847 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 848 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 849 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 850 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 851 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 852 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 853 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 854 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 855 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 856 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 857 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 858 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 859 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 860 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 861 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 862 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 863 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 864 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 865 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 866 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 867 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 868 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 869 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 870 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 871 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 872 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 873 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 874 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 875 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 876 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 877 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 878 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 879 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 880 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 881 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 882 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 883 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 884 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 885 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 886 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 887 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 888 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 889 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 890 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 891 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 892 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 893 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 894 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 895 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 896 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 897 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 898 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 899 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 900 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 901 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 902 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 903 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 904 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 905 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 906 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 907 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 908 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 909 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 910 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 911 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 912 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 913 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 914 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 915 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 916 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 917 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 918 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 919 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 920 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 921 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 922 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 923 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 924 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 925 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 926 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 927 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
instance Random 928 where
  mkRandomN = mkAutoStepLFSR ∘ mkLFSRRandSeedN
