typedef union tagged {
   union tagged {
      Bool First;
      void Second;
   } OneTwo;
   void Three;
} TaggedUnionTagged;

