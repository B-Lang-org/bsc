function Action f();
  action
    x = 3;
  endaction
endfunction
