`define is 1
`define fs 500
`define full sysFromReal_1_500

`include "FromReal.bsv"
