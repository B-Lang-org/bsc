import Sub2::*;

interface Ifc1;
   (* prefix="" *)
   interface Ifc2 wr;
endinterface

