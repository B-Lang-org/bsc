function bit[3:0] f();
  bit[3:0] x = 3, y, z = 5;
  y = 4;
  f = x + y + z;
endfunction
