(* synthesize *)
module sysInvalid_Int_Oct ();
   Reg#(Bit#(4)) rg <- mkReg('o777);
endmodule
