
(* synthesize, synthesize *)
module sysMultipleSameAttribModule();
endmodule
