// Bug 681

module mkModIfc_TooFewArgs_TopLevel(Reg);
endmodule
