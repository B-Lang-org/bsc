import Vector::*;

(* synthesize *)
(* gate_input_clocks="clks" *)
module sysGateInputClocks_VecClock ( Vector#(2,Clock) clks,
                                     Empty ifc );
endmodule

