package CircTop;

import CircPkg::*;

export CircPkg::*;

endpackage

