
interface Ifc;
 method Action check ((* port="y " *)Bool x);
endinterface

