
typedef List#(A) A;

