
(* synthesized *)
module sysT1();
endmodule

