ActionValue#(Bool) av;
av =
  actionvalue
    bit[3:0] x = 3;
    return True;
  endactionvalue;

