package EmptyCase() where

x :: Bool
x = True

emptyCase :: Bool
emptyCase = case x of {};