package UTF8Cons1(Ptak(..)) where

data Ptak = Żuraw | Gżegżółka | Gołąb

