Bit#(8) x = 5;