package UTF8MultilineComment(foo) where

{-
   comment ·
   with · a · non-ASCII
   · symbol
   zażółć gęsią jaźń
   ここには何でも書いていい
 -}

foo :: (Bits a sza) => a -> a
foo = unpack `compose` pack

