package OneArgMissingOne () where

x :: Bit
x = _

