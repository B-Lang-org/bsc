module sysExplictBool();
   Bool x=99;
   Bool y=10;
endmodule
