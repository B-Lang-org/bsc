package ClassDefParamGivenNonNumUsedNum () where

class (Foo :: * -> *) a where
    bar :: Bit a

