package TypeAliasParamGivenNumUsedNonNum () where

data (Foo :: * -> *) a = Bar a

type (Baz :: # -> *) b = Foo b

