-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EUnknownSize.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the EUnknownSize error of the bluespec
-- compiler (Bit Vector of unknown size introduced near this location)
--
-----------------------------------------------------------------------



package EUnknownSize2 () where

x :: Bit n
x = if x==0 then 1 else 0





