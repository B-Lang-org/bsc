(* synthesize *)
module sysPrintType();

  Bool b = True;
  messageM(printType(typeOf(b)));

endmodule

