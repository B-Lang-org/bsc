package DanglingDecimal where

x :: Integer
x = 0.
