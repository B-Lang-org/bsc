package Fake_WFilePackageNameMismatch_Sub(foo) where

foo :: Integer
foo = 1
