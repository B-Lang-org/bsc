package Bug353_Type where

data Foo a b = Foo b
