package Export(_) where

