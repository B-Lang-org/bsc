function Bit#(1) f();
   Bit#(TSub#(3,4)) x = 0;
   return x;
endfunction

