// Comment

`line(/file/path,4,1 1,0)

Bool b = True;
