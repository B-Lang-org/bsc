(* clock_prefix="" *)
module sysEmptyCLKAttrib ();
endmodule

