package BindDummyLambda () where

x :: Bool -> Int 32
x = \_ -> _

