package RecDeriveDataOneArgManyTypeArgs () where

data Foo a = F (Foo a) deriving (Eq)

