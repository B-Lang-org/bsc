(* synthesize *)
module sysInputArg_Unused #(Bit#(16) b) ();
endmodule

