package Empty () where

interface Null = {}

mkEmpty :: Module Null
mkEmpty =
    module
