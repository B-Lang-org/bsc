package 風呂敷;

endpackage: 風呂敷
