(* synthesize *)
module sysPropDeduce_NoUse ();
endmodule

