// Accellera Standard V2.8.1 Open Verification Library (OVL).
// Accellera Copyright (c) 2005-2014. All rights reserved.

`include "std_ovl_defines.h"

`module ovl_frame (clock, reset, enable, start_event, test_expr, fire);

  parameter severity_level      = `OVL_SEVERITY_DEFAULT;
  parameter min_cks             = 0;
  parameter max_cks             = 0;
  parameter action_on_new_start = `OVL_ACTION_ON_NEW_START_DEFAULT;
  parameter property_type       = `OVL_PROPERTY_DEFAULT;
  parameter msg                 = `OVL_MSG_DEFAULT;
  parameter coverage_level      = `OVL_COVER_DEFAULT;

  parameter clock_edge     = `OVL_CLOCK_EDGE_DEFAULT;
  parameter reset_polarity = `OVL_RESET_POLARITY_DEFAULT;
  parameter gating_type    = `OVL_GATING_TYPE_DEFAULT;

  input                          clock, reset, enable;
  input                          start_event;
  input                          test_expr;
  output [`OVL_FIRE_WIDTH-1:0]   fire;

  // Parameters that should not be edited
  parameter assert_name = "OVL_FRAME";

  `include "std_ovl_reset.h"
  `include "std_ovl_clock.h"
  `include "std_ovl_cover.h"
  `include "std_ovl_task.h"
  `include "std_ovl_init.h"

`ifdef OVL_SYNTHESIS
`else
  // Sanity Checks
  initial begin
    if (~((action_on_new_start == `OVL_IGNORE_NEW_START)   ||
          (action_on_new_start == `OVL_RESET_ON_NEW_START) ||
          (action_on_new_start == `OVL_ERROR_ON_NEW_START)))
    begin
      ovl_error_t(`OVL_FIRE_2STATE,"Illegal value set for parameter action_on_new_start");
    end
    //
    if ((max_cks > 0) && (min_cks > max_cks)) begin
       ovl_error_t(`OVL_FIRE_2STATE,"Illegal parameter values set where min_cks > max_cks");
    end
  end
`endif

`ifdef OVL_VERILOG
  `include "./vlog95/assert_frame_logic.v"
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.3
`endif

`ifdef OVL_SVA
  `include "./sva05/assert_frame_logic.sv"
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.3
`endif

`ifdef OVL_PSL
  assign fire = {`OVL_FIRE_WIDTH{1'b0}}; // Tied low in V2.3
  `include "./psl05/assert_frame_psl_logic.v"
`else
  `endmodule // ovl_frame
`endif
