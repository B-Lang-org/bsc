package IfLiftingTwoArg(sysIfLiftingTwoArg) where

-- Lifting of if-branches: `b.set False' and `b.set True' on two sides
-- of the `if' should be lifted out to `b.set (nosplitIf a False True)'

import RegFile 

sysIfLiftingTwoArg :: Module Empty
sysIfLiftingTwoArg =
  module
    a :: Reg Bool
    a <- mkRegU
    b :: RegFile (Bit 5) (Int 32) <- mkRegFileFull
    rules
        when True ==> if a then b.upd 9 17 else b.upd 12 19

