module mkModIfc_TooFewArgs_Local();
   module mkMod(Reg); endmodule
endmodule
