package IfcArgNamesUpper where

interface Foo =
    foo :: Bool -> Action {-# arg_names = [FOOBAR] #-}

{-# synthesize mkFoo #-}
mkFoo :: Module Foo
mkFoo = return _
