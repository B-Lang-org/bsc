
(* synthesize *)
module sysLiteral_TooLarge();
   Reg#(Bit#(11)) rg <- mkReg('h800);
endmodule

