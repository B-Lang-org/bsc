import Basic::*;
export Basic::*;

