`include <defines1

Bool x = message(`V, True);

