package TypeAliasResGivenNumIsNonNumParam () where

type (Foo :: * -> #) a = a

