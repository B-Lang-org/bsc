import MyRAM::*;

(* synthesize *)
module mkTest (MyRAM#(Bit#(8),Bit#(16)));
   return ?;
endmodule

