// These comments should not be lost

`define y endmodule

`define m(x) x

module sysTest();

`m(`y)

// more here