(* synthesize *)
module sysDigitToInteger_Bad();
   rule r;
      $display(digitToInteger("a"));
   endrule
endmodule
