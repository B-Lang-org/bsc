typedef "Foo" Name;

function Bool isName (String x);
   return (Name == x);
endfunction
