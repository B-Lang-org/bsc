// Valid attribute is wrong place

(* synthesize *)
interface Foo ;
   method Action start () ;
endinterface 
      
module sysT2();
endmodule

