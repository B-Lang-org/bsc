package DegreePrimeVar2() where

a´ :: a -> a
a´ = id
