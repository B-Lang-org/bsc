module sysActions();
   rule test1;
      False;
   endrule
   rule test2;
      True;
   endrule
endmodule
