module mkProvisoBaseMismatch_Local();
   module mkMod(Reg#(t))
      provisos(Add#(1,j,t));
   endmodule
endmodule
