typedef union tagged {
   Bool First;
   void First;
   void Second;
} TaggedUnionSimple;

