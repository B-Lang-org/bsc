typedef union tagged {
  a T1;
  b T2;
} U #(type a, type b, type a);

