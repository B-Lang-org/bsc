package TestExcludeBad where

import Exclude

d :: Integer
d = b + a * b