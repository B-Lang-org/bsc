(* synthesize *)
module mkAbstractDerivePosition();
   primError(?, "this is an error message");
endmodule
