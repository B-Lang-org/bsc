-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EBigLiteral.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the EBigLiteral error of the bluespec
-- compiler (Literal {literal} does not fit in # bits)
--
-- Generates error if code is requested for mkGCD
-----------------------------------------------------------------------



package EBigLiteral (GCD(..), mkGCD) where

-- import UInt

interface GCD =
    start  :: UInt 2 -> UInt 2 -> Action
    result :: UInt 2

mkGCD :: Module GCD
mkGCD =
    module
        x :: Reg (UInt 2)
        x <- mkRegU

        y :: Reg (UInt 2)
        y <- mkReg 5

        rules
          "Swap":
            when x > y, y /= 0
              ==> action
                      x := y
                      y := x

          "Subtract":
            when x <= y, y /= 0
              ==> action
                      y := y - x

        interface
            start ix iy = action
                              x := ix
                              y := iy
                          when y == 0
            result = x when y == 0


