`define comment //
`comment
