
import "BDPI" my_C_or = function Bit#(8) my_or (Bit#(8) x, Bit#(8) y);

