interface Foo#(numeric type a);
endinterface

module mkInterfacePartialKind(Foo#(1));
endmodule

