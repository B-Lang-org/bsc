/*
 * any unicode is ok in comments
 *
 * comment
 * · with · a · non-ASCII
 * · symbol
 * zażółć gęsią jaźń
 * ここには何でも書いていい
 */

export foo;

function a foo(a x);
    return x;
endfunction: foo

