
interface Ifc;
 method Action check ((* port="" *)Bool x);
endinterface

