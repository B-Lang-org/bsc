module sysAmbigTCon_TDiv (Reg#(Bit#(TDiv#(x,y))));
endmodule
