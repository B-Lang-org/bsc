
`define m(x
) x

Bool b = `m(True);

Bool b2 = `m(False);
