export Cvijet;

// uppercase and titlecase lj digraphs can start constructors

typedef union tagged {
   Bool ǇIǇAN;
   void  ǈiǉan;
} Cvijet;

