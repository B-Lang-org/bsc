module ThreeClocks(CLK_a, CLK_b, CLK_c);

   output CLK_a;
   output CLK_b;
   output CLK_c;

   wire CLK_a = 0;
   wire CLK_b = 0;
   wire CLK_c = 0;
   
endmodule // ThreeClocks
