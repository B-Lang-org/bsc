Bool x = True | True;

