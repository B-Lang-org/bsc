
module Empty(CLK, RST_N);
   input     CLK;
   input     RST_N;


endmodule

