package NumPlusOne () where

x :: 1 Bool
x = _

