import Vector::*;

// Test that we don't get two messages about "replicateM"
export Vector::*;
export replicateM;
export replicateM;

