module sysAmbigTCon_TExp (Reg#(Bit#(TExp#(n))));
endmodule
