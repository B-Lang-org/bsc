function bit[3:0] f();
  bit[3:0] x;
  x = x;
  f = x;
endfunction
