package DegreePrimeVar4(a´) where

a´ :: a -> a
a´ = id
