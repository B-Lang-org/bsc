import ClassWithDefault_Interface::*;

module sysImportClassWithDefault_Interface (Reg#(Bit#(8)));
   Reg#(Bit#(8)) x <- cmod;
   return x;
endmodule
