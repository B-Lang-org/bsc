package Undet1(sysUndet1) where

sysUndet1 :: Module Empty
sysUndet1 =
  module
    x :: Reg (Bit 27) <- mkReg 2
    counter :: Reg (Bit 16) <- mkReg 0

    rules 
      when True ==> counter := counter + 1
      when True ==> if (counter < 16) then displayHex(x :: Bit 27) else $finish 0
      when (counter == 4) ==> x := _
      when (counter == 8) ==> x := 5
