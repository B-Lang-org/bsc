package DupObj;

Bool x = False;

endpackage
