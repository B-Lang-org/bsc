Cpreprocess.bsv