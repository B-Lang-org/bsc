module mkFoo();
  rule bogus1;
  endrule
endmodule
