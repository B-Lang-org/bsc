Integer foo;
foo = -5;
