package Overlap1(sysOverlap1) where

class Displayable a where
   display :: a -> Action

instance (Bits a sa) => Displayable a 
   where
     display a = $display "Bits %h" a

instance (Displayable a) => Displayable (Maybe a)
   where 
     display (Valid a) = action
                           $write "Valid "
                           display a
     display (Invalid) = $display "Invalid"

{-# verilog sysOverlap1 #-}
sysOverlap1 :: Module Empty
sysOverlap1 = 
  module
    x :: Reg (Maybe (Bit 17)) <- mkReg Invalid
    rules
      "test":
         when True  ==>
           action
               display x
               $finish 0
