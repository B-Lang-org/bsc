package RecDeriveDataInsideList () where

data Foo = F (List Foo) deriving (Eq)

