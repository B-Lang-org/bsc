module sysExplictRules();
   Rules r=rules rule test; noAction; endrule endrules;
   Rules a=True;
   Rules b=False;
endmodule
