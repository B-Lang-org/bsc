package UndefinedTask() where

foo :: Action
foo = $foobar 17