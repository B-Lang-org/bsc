`define FOO

`ifdef

FOO
Bool x = True;
`endif

