
import Basic::*;

export Basic::*;

function Bool myFn1(Integer x);
  return (x > 2);
endfunction

typedef enum { A, B } S;

