module mkTest ();
  Tuple3#(Bool, Integer, Bit#(8)) { .* , .* , .* } = tuple3(True,1,2);
endmodule
