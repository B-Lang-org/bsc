(* synthesize *)
module sysInitialBlocks();
    Reg#(int) r <- mkRegU();
endmodule
