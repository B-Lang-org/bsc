
interface Ifc;
 (* ready = "always" *)
 method Bool check ();
endinterface

(* synthesize *)
module mkKeyword (Ifc);
endmodule
