package LexPos where

x :: Integer
x = 5 + 9 + "foo"

y :: Integer
y = 0x5 + 0xA + "bar"