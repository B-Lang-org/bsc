/////////////////////////////////////////////////////////////////////////
/* Defines all the constants related to this module
*/

package Defines;

  // Aspect ratio info
  Bit#(4)  eXTENDED_PAR = 4'b1111;


  // Video object layer shape
  Bit#(2)  rECTANGULAR  = 2'b00 ;
  Bit#(2)  bINARY       = 2'b01 ;
  Bit#(2)  bINARY_ONLY  = 2'b10 ;
  Bit#(2)  gRAYSCALE    = 2'b11 ;

  Bit#(2)  sTATIC       = 2'b01 ;
  Bit#(2)  gMC          = 2'b10 ;


  Bit#(2)  aUX_COMP_COUNT  = 2'b01 ;
  
typedef enum {IDLE,START,WAIT,SUSPEND } PSstates
          deriving (Eq,Bits);  

typedef enum {EXTENDED_PAR} AspectRatioStates
          deriving (Eq,Bits);  

typedef enum {NOTUSED,TYPE1,TYPE2,TYPE3,TYPE4} FLC_type
          deriving (Eq,Bits);  

typedef enum {IDLE,
              SUSPEND,
              RESUME,
              VIDEO_OBJECT_LAYER0,
			  VIDEO_OBJECT_LAYER1,
			  VIDEO_OBJECT_LAYER1_1,
			  VIDEO_OBJECT_LAYER1_2,
			  VIDEO_OBJECT_LAYER2,
			  VIDEO_OBJECT_LAYER2_0,
			  VIDEO_OBJECT_LAYER2_1,
			  VIDEO_OBJECT_LAYER2_1_0,
			  VIDEO_OBJECT_LAYER3,
			  VIDEO_OBJECT_LAYER3_0,
			  VIDEO_OBJECT_LAYER3_0_1,
			  VIDEO_OBJECT_LAYER3_0_2,
			  VIDEO_OBJECT_LAYER3_1,
			  VIDEO_OBJECT_LAYER3_2,
			  VIDEO_OBJECT_LAYER4,
			  VIDEO_OBJECT_LAYER4_0_1,
			  VIDEO_OBJECT_LAYER4_1,
			  VIDEO_OBJECT_LAYER4_1_1,
			  VIDEO_OBJECT_LAYER4_1_2,
			  VIDEO_OBJECT_LAYER4_1_3,
			  VIDEO_OBJECT_LAYER4_2,
			  VIDEO_OBJECT_LAYER4_2_1,
			  VIDEO_OBJECT_LAYER5_0_1,
			  VIDEO_OBJECT_LAYER5_1,
			  VIDEO_OBJECT_LAYER5_1_1,
			  VIDEO_OBJECT_LAYER5_1_1_1,
			  VIDEO_OBJECT_LAYER5_1_2,
			  VIDEO_OBJECT_LAYER5_1_2_1,
			  VIDEO_OBJECT_LAYER5_1_3,
			  VIDEO_OBJECT_LAYER5_1_4,
			  VIDEO_OBJECT_LAYER5_1_5,
			  VIDEO_OBJECT_LAYER5_1_6,
			  VIDEO_OBJECT_LAYER5_1_7,
			  VIDEO_OBJECT_LAYER5_1_8,
			  VIDEO_OBJECT_LAYER5_1_9,
			  VIDEO_OBJECT_LAYER5_1_10,
			  VIDEO_OBJECT_LAYER5_1_11,
			  VIDEO_OBJECT_LAYER5_2,
			  VIDEO_OBJECT_LAYER5_2_1,
			  VIDEO_OBJECT_LAYER5_2_2,
			  VIDEO_OBJECT_LAYER5_2_2_0,
			  VIDEO_OBJECT_LAYER5_3,
			  VIDEO_OBJECT_LAYER5_3_1,
			  VIDEO_OBJECT_LAYER5_4,
			  VIDEO_OBJECT_LAYER5_4_1,
			  VIDEO_OBJECT_LAYER5_5,
			  VIDEO_OBJECT_LAYER5_5_1,
			  VIDEO_OBJECT_LAYER5_6,
			  VIDEO_OBJECT_LAYER5_6_0,
			  VIDEO_OBJECT_LAYER5_6_1,
			  VIDEO_OBJECT_LAYER5_6_2,
			  VIDEO_OBJECT_LAYER5_6_1_1,
			  VIDEO_OBJECT_LAYER6,
			  VIDEO_OBJECT_LAYER7,
			  VIDEO_OBJECT_LAYER9,
			  VIDEO_OBJECT_LAYER9_1_0,
			  VIDEO_OBJECT_LAYER9_2,
			  VIDEO_OBJECT_LAYER9_2_0,
			  VIDEO_OBJECT_LAYER9_3,
			  VIDEO_OBJECT_LAYER9_3_1,
			  VIDEO_OBJECT_LAYER9_4,
			  VIDEO_OBJECT_LAYER9_4_1,
			  VIDEO_OBJECT_LAYER9_5,
			  VIDEO_OBJECT_LAYER9_5_0,
			  VIDEO_OBJECT_LAYER10,
			  VIDEO_OBJECT_LAYER10_1_0,
			  VIDEO_OBJECT_LAYER10_2,
			  VIDEO_OBJECT_LAYER10_2_0,
			  VIDEO_OBJECT_LAYER10_3,
			  VIDEO_OBJECT_LAYER10_3_0,
			  VIDEO_OBJECT_LAYER11,
			  VIDEO_OBJECT_LAYER11_1,
			  VIDEO_OBJECT_LAYER11_1_0,
			  VIDEO_OBJECT_LAYER11_2,
			  VIDEO_OBJECT_LAYER11_2_0,
			  VIDEO_OBJECT_LAYER11_3,
			  VIDEO_OBJECT_LAYER11_4,
			  VIDEO_OBJECT_LAYER11_5,
			  VIDEO_OBJECT_LAYER11_6,
			  VIDEO_OBJECT_LAYER11_7,
			  VIDEO_OBJECT_LAYER12,
			  VIDEO_OBJECT_LAYER12_1_0,
			  VIDEO_OBJECT_LAYER12_2,
			  VIDEO_OBJECT_LAYER12_2_0,
			  VIDEO_OBJECT_LAYER12_3,
			  VIDEO_OBJECT_LAYER12_3_0,
			  VIDEO_OBJECT_LAYER13,
			  VIDEO_OBJECT_LAYER13_1,
			  VIDEO_OBJECT_LAYER13_1_0,
			  VIDEO_OBJECT_LAYER14,
			  VIDEO_OBJECT_LAYER14_1_0,
			  VIDEO_OBJECT_LAYER15,
			  VIDEO_OBJECT_LAYER15_1_0,
			  VIDEO_OBJECT_LAYER16,
			  VIDEO_OBJECT_LAYER17,
			  VIDEO_OBJECT_LAYER17_1_0,
			  VIDEO_OBJECT_LAYER18,
			  VIDEO_OBJECT_LAYER18_1_0,
			  VIDEO_OBJECT_LAYER19,
			  VIDEO_OBJECT_LAYER19_1_0,
			  VIDEO_OBJECT_LAYER19_2,
			  VIDEO_OBJECT_LAYER19_2_0,
			  VIDEO_OBJECT_LAYER20,
			  VIDEO_OBJECT_LAYER20_1_0,
			  VIDEO_OBJECT_LAYER20_2,
			  VIDEO_OBJECT_LAYER20_2_0,
			  VIDEO_OBJECT_LAYER21,
			  VIDEO_OBJECT_LAYER21_1_0,
			  VIDEO_OBJECT_LAYER21_1,
			  VIDEO_OBJECT_LAYER22,
			  VIDEO_OBJECT_LAYER22_1_0,
			  VIDEO_OBJECT_LAYER23,
			  VIDEO_OBJECT_LAYER24_1_0,
			  VIDEO_OBJECT_LAYER24,
			  VIDEO_OBJECT_LAYER24_2,
			  VIDEO_OBJECT_LAYER25,
			  VIDEO_OBJECT_LAYER25_1,
			  VIDEO_OBJECT_LAYER25_1_1,
			  VIDEO_OBJECT_LAYER26,
			  VIDEO_OBJECT_LAYER26_1_1,
			  VIDEO_OBJECT_LAYER27,
			  VIDEO_OBJECT_LAYER27_1_1,
			  VIDEO_OBJECT_LAYER28,
			  VIDEO_OBJECT_LAYER28_1_1,
			  VIDEO_OBJECT_LAYER29,
			  VIDEO_OBJECT_LAYER29_1_1,
			  VIDEO_OBJECT_LAYER30,
			  VIDEO_OBJECT_LAYER30_1,
			  VIDEO_OBJECT_LAYER30_1_1,
			  VIDEO_OBJECT_LAYER31_1,
			  VIDEO_OBJECT_LAYER31_1_1,
			  VIDEO_OBJECT_LAYER31_2,
			  VIDEO_OBJECT_LAYER31_2_1,
			  VIDEO_OBJECT_LAYER32,
			  VIDEO_OBJECT_LAYER32_2,
			  VIDEO_OBJECT_LAYER32_1_1,
			  VIDEO_OBJECT_LAYER32_2_1,
			  VIDEO_OBJECT_LAYER32_3,
			  VIDEO_OBJECT_LAYER32_3_1,
			  VIDEO_OBJECT_LAYER32_4,
			  VIDEO_OBJECT_LAYER32_5,
			  VIDEO_OBJECT_LAYER32_6,
			  VIDEO_OBJECT_LAYER32_6_1,
			  VIDEO_OBJECT_LAYER33,
			  VIDEO_OBJECT_LAYER33_1_1,
			  VIDEO_OBJECT_LAYER33_1_2,
			  VIDEO_OBJECT_LAYER33_2_1,
			  VIDEO_OBJECT_LAYER33_2,
			  VIDEO_OBJECT_LAYER33_3,
			  VIDEO_OBJECT_LAYER33_4,
			  VIDEO_OBJECT_LAYER34,
			  VIDEO_OBJECT_LAYER34_1,
			  VIDEO_OBJECT_LAYER34_1_1,
			  VIDEO_OBJECT_LAYER34_2,
			  VIDEO_OBJECT_LAYER34_2_1,
			  VIDEO_OBJECT_LAYER34_3,
			  VIDEO_OBJECT_LAYER34_4,
			  VIDEO_OBJECT_LAYER35,
			  VIDEO_OBJECT_LAYER35_1,
			  VIDEO_OBJECT_LAYER36,
			  VIDEO_OBJECT_LAYER37,
			  VIDEO_OBJECT_LAYER37_1,
			  VIDEO_OBJECT_LAYER37_1_0,
			  VOL_NEXT_START_CODE_DET,
			  USER_DATA,
			  USER_DATA1,
			  GROUP_OF_VOP,
			  GROUP_OF_VOP_1,
			  GROUP_OF_VOP_1_0,
			  GROUP_OF_VOP_2,
			  GROUP_OF_VOP_2_0,
			  GROUP_OF_VOP_3,
			  GROUP_OF_VOP_3_0,
			  GROUP_OF_VOP_4,
			  GROUP_OF_VOP_5,
			  GROUP_OF_VOP_5_0,
			  GROUP_OF_VOP_5_1_0,
			  GROUP_OF_VOP_5_1,
			  VOP_STATE,
			  VOP_STATE_0,
			  VOP_STATE_0_1,
			  VOP_STATE_1,
			  VOP_STATE_1_0,
			  VOP_STATE_2,
			  VOP_STATE_CAL_FVTI,
			  VOP_STATE_2_0,
			  VOP_STATE_2_1,
			  VOP_STATE_2_1_0,
			  VOP_STATE_2_2,
			  VOP_STATE_2_3,
			  VOP_STATE_2_4,
			  VOP_STATE_2_4_0,
			  VOP_STATE_3,
			  VOP_STATE_3_0,
			  VOP_STATE_3_0_0,
			  VOP_STATE_3_1,
			  VOP_STATE_3_1_0,
			  VOP_STATE_4,
			  VOP_STATE_4_0,
			  VOP_STATE_4_0_0,
			  VOP_STATE_5,
			  VOP_STATE_5_1,
			  VOP_STATE_4_READ_VOP_COMPLEXITY_ESTIMATION_HEADER,
			  VOP_STATE_6,
			  VOP_STATE_6_0,
			  VOP_STATE_7,
			  VOP_STATE_8,
			  VOP_STATE_8_0,
			  VOP_STATE_9,
			  VOP_STATE_10,
			  VOP_STATE_10_0,
			  VOP_STATE_11,
			  VOP_START_CODE_DET,
			  DATA_PARTITIONED_MST,
			  COMBINED_MST0,
			  COMBINED_MST_0_1,
			  COMBINED_MST_0_2,
			  COMBINED_MST,
			  MB_not_coded_wait_state,
			  MB_not_coded_wait_state_1,
			  MB_not_coded_wait_state_2,
			  WAIT64,
			  JUST_WAIT64,
			  MB_STATE_1,
			  MB_STATE_1_0,
			  MB_STATE_2,
			  MB_STATE_3,
			  MB_STATE_3_0,
			  MB_STATE_4,
			  MB_STATE_5,
			  MB_STATE_5_0,
			  MB_STATE_6,
			  MB_STATE_7,
			  MB_STATE_7_0,
			  MB_STATE_8,
			  MB_STATE_9,
			  MB_STATE_9_0,
			  MB_STATE_10,
			  MST_STATE_0,
			  MV_STATE_1,
			  MV_STATE_2,
			  MV_STATE_2_0,
			  MV_STATE_2_1,
			  MV_STATE_2_1_0,
			  MV_STATE_2_2,
			  MV_STATE_2_2_0,
			  MV_STATE_3,
			  MV_STATE_4,
			  MV_STATE_4_0,
			  MV_STATE_5,
			  MV_STATE_6,
			  MV_STATE_6_0,
			  MV_STATE_6_1,
			  MV_STATE_6_1_0,
			  MV_STATE_6_2,
			  MV_STATE_6_2_0,
			  MV_STATE_7,
			  MV_STATE_8,
			  MV_STATE_8_0,
			  MV_STATE_10,
			  EXEC_MV_PREDICTION,
			  EXEC_MV_PREDICTION1,
			  EXEC_4MV_PREDICTION,
			  EXEC_4MV_PREDICTION1,
			  EXEC_4MV_PREDICTION2,
			  EXEC_4MV_PREDICTION3,
			  UPDATE_MV_BUFFER,
			  MB_BLK_STATE,
			  MB_BLK_STATE_0,
			  MB_BLK_STATE_00,
			  MB_BLK_STATE_00_0,
			  MB_BLK_STATE_1,
			  MB_BLK_STATE_1_0,
			  MB_BLK_STATE_2,
			  MB_BLK_STATE_2_0,
			  MB_BLK_STATE_2_1,
			  MB_BLK_STATE_2_1_0,
			  MB_BLK_STATE_3,
			  MB_BLK_STATE_4,
			  MB_BLK_STATE_4_0,
			  MB_BLK_STATE_5,
			  MB_BLK_STATE_6,
			  MB_BLK_STATE_6_0,
			  MB_BLK_STATE_7,
			  MB_BLK_STATE_7_0,
			  MB_BLK_STATE_7_1,
			  MB_BLK_STATE_7_1_0,
			  MB_BLK_STATE_8,
			  MB_BLK_STATE_9,
			  MB_BLK_STATE_9_0,
			  MB_BLK_STATE_10,
			  MB_BLK_STATE_11,
			  MB_BLK_STATE_11_0,
			  MB_BLK_STATE_12,
			  MB_BLK_STATE_DCTVlc,
			  MB_BLK_STATE_DCTVlc_0,
			  MB_BLK_STATE_DCTVlc_0_0,
			  DecodeVLCIntraTable1,
			  DecodeVLCIntraTable2,
			  DecodeVLCIntraTable3,
			  DecodeVLCIntraTable4,
			  DecodeVLCIntraTable5,
			  DecodeVLCIntraTable6,
			  DecodeVLCIntraTable7,
			  DecodeVLCIntraTable8,
			  DecodeVLCIntraTable9,
			  DecodeVLCInterTable1,
			  DecodeVLCInterTable2,
			  DecodeVLCInterTable3,
			  DecodeVLCInterTable4,
			  DecodeVLCInterTable5,
			  DecodeVLCInterTable6,
			  DecodeVLCInterTable7,
			  DecodeVLCInterTable8,
			  DecodeVLCInterTable9,
			  Fixed_length_code,
			  MB_BLK_STATE_FLC_Type3,
			  MB_BLK_STATE_FLC_Type3_0,
			  MB_BLK_STATE_FLC_Type3_1,
			  MB_BLK_STATE_FLC_Type3_1_0,
			  MB_BLK_STATE_FLC_Type3_2,
			  MB_BLK_STATE_FLC_Type3_2_0,
			  EXEC_ACDC_PREDICTION,
			  EXEC_ACDC_PREDICTION_INTER,
			  EXEC_ACDC_PREDICTION1,
			  EXEC_ACDC_PREDICTION2,
			  EXEC_ACDC_PREDICTION3,
			  CHECK_RESYNC_MARKER,
			  CHECK_RESYNC_MARKER0,
			  CHECK_RESYNC_MARKER0_0,
			  CHECK_RESYNC_MARKER0_1,
			  CHECK_RESYNC_MARKER0_1_0,
			  CHECK_RESYNC_MARKER_0,
			  CHECK_RESYNC_MARKER1,
			  CHECK_RESYNC_MARKER2,
			  CHECK_RESYNC_MARKER2_0,
			  CHECK_RESYNC_MARKER3,
			  VIDEO_PACKET_HEADER,
			  VIDEO_PACKET_HEADER0,
			  VIDEO_PACKET_HEADER_1_0,
			  VIDEO_PACKET_HEADER_1,
			  VIDEO_PACKET_HEADER_2_0,
			  VIDEO_PACKET_HEADER_2,
			  START_CODE_DET,
			  START_CODE_DET0,
			  START_CODE_DET_1,
			  START_CODE_DET_1_0
			  } VideoSt
          deriving (Eq,Bits); 

typedef Tuple2#(Bit#(8), Bit#(8)) DtSrct ;

typedef Tuple7#(Bit#(9),Bit#(1),Bit#(4),Bit#(2),Bit#(1),Bit#(48),Bit#(48)) Mbheadertype;
typedef Tuple6#(Bit#(12),Bit#(12),Bit#(12),Bit#(12),Bit#(12),Bit#(12)) MVtype;

endpackage : Defines
