int someint;
someint = 1;

Int#(16) otherint;
otherint = someint;
