function t3 fn(t1 v, t2 v);
  return ?;
endfunction
