module mkTest();
  Reg#(Bit#(6)) r;
  mkReg#(y) the_r;
endmodule
