import ReExportItems_Q::*;

// test that the type made it
AB b2 = B;

// test that the variable made it
Bool aOK = a == A;


