export 鳥;

// kanji are not unicode uppercase letters

typedef union tagged {
   Bool 鶴;
   void 梟;
} 鳥;

