Integer x = 'h5xx7;
