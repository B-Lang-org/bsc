package Expr_Where () where

x :: Bool
x = _ where v = True

