package NoType where

x = 5