module test1 ();
   Bool f = 13;
endmodule
