// polymorphic function definition

function a id(a thing);
  id = thing;
endfunction
