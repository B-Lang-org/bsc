typeclass C#(numeric type a, type b);
   function Bit#(a) cf();
   function b f2(b x);
endtypeclass

