`include "DupInclude.defines"

Bool y = x;

