module mkTest1 (Empty);
    Reg#(Int#(32)) x();
    mkReg#(?,?) the_x(x);
endmodule
