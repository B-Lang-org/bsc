interface Ifc;
endinterface

module sysBug547(Ifc);
  rule bogus;
  endrule
endmodule
