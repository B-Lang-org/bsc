package Types_NonNamed where

-- BSC represents this as a constructor of one argument
-- that is a struct with fields named "_1" and "_2".
-- However, this should not be visible to users.
--
data Foo = Bar Bool Bool
