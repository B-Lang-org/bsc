package InstanceSplit where

import Vector
import BuildVector
import SplitPorts
import CShow

struct Foo =
  x :: Int 8
  y :: Int 8
 deriving (Bits)

instance SplitPorts Foo (Port (Int 8), Port Bool, Port (Bit 7)) where
  splitPorts x = (Port x.x, Port (x.y > 0), Port $ truncate $ pack x.y)
  unsplitPorts (Port x, Port s, Port y) = Foo { x = x; y = (if s then id else negate) $ unpack $ zeroExtend y; }
  portNames _ base = Cons (base +++ "_x") $ Cons (base +++ "_ysign") $ Cons (base +++ "_yvalue") Nil

struct Bar =
  v :: Vector 3 Bool
  w :: (Bool, UInt 16)
  z :: Foo
 deriving (Bits)

-- XXX would be nice to be able to derive this
instance (ShallowSplitPorts Bar p) => SplitPorts Bar p where
  splitPorts = shallowSplitPorts
  unsplitPorts = shallowUnsplitPorts
  portNames = shallowSplitPortNames

struct Baz =
  a :: Maybe Foo
  b :: Bar
  c :: Vector 3 (Vector 8 Foo, Bar)
  d :: ()
  e :: Vector 0 Foo
 -- No Bits instance needed

-- XXX would be nice to be able to derive this
instance (ShallowSplitPorts Baz p) => SplitPorts Baz p where
  splitPorts = shallowSplitPorts
  unsplitPorts = shallowUnsplitPorts
  portNames = shallowSplitPortNames

interface SplitTest =
  putFoo :: Foo -> Action
  putBar :: Bar -> Action {-# prefix = "PUT_BAR" #-}
  putFooBar :: Foo -> Bar -> Action {-# arg_names = ["fooIn", "barIn"] #-}
  putFoos :: (Vector 50 Foo) -> Action
  putBaz :: Baz -> Action


{-# synthesize mkInstanceSplitTest #-}
mkInstanceSplitTest :: Module SplitTest
mkInstanceSplitTest =
  module
    interface
      putFoo x = $display "putFoo: " (cshow x)
      putBar x = $display "putBar: " (cshow x)
      putFooBar x y = $display "putFooBar: " (cshow x) " " (cshow y)
      putFoos x = $display "putFoos: " (cshow x)
      putBaz x = $display "putBaz: " (cshow x)

{-# synthesize sysInstanceSplit #-}
sysInstanceSplit :: Module Empty
sysInstanceSplit =
  module
    s <- mkInstanceSplitTest
    i :: Reg (UInt 8) <- mkReg 0
    rules
      when True ==> i := i + 1
      when i == 0 ==> s.putFoo $ Foo { x = 1; y = 2; }
      when i == 1 ==> s.putBar $ Bar { v = vec True False True; w = (True, 0x1234); z = Foo { x = 3; y = 4; } }
      when i == 2 ==> s.putFooBar (Foo { x = 5; y = 6; }) (Bar { v = vec False True False; w = (False, 0x5678); z = Foo { x = 7; y = 8; } })
      when i == 3 ==> s.putFoos $ genWith $ \ j -> Foo { x = fromInteger $ 9 + j / 2; y = fromInteger $ 10 - 2*j / 3; }
      when i == 4 ==> s.putBaz $ Baz { a = Just $ Foo { x = 9; y = 10; }; b = Bar { v = vec True False False; w = (True, 0x1234); z = Foo { x = 3; y = 4; }; }; c = vec (vec (Foo { x = 11; y = 12; }) (Foo { x = 13; y = 14; }) (Foo { x = 15; y = 16; }) (Foo { x = 17; y = 18; }) (Foo { x = 19; y = 20; }) (Foo { x = 21; y = 22; }) (Foo { x = 23; y = 24; }) (Foo { x = 25; y = 26; }), Bar { v = vec True False True; w = (True, 0xBEEF); z = Foo { x = 3; y = 4; } }) (vec (Foo { x = 27; y = 28; }) (Foo { x = 29; y = 30; }) (Foo { x = 31; y = 32; }) (Foo { x = 33; y = 34; }) (Foo { x = 35; y = 36; }) (Foo { x = 37; y = 38; }) (Foo { x = 39; y = 40; }) (Foo { x = 41; y = 42; }), Bar { v = vec True False True; w = (True, 0x4321); z = Foo { x = 123; y = 42; } }) (vec (Foo { x = 43; y = 44; }) (Foo { x = 45; y = 46; }) (Foo { x = 47; y = 48; }) (Foo { x = 49; y = 50; }) (Foo { x = 51; y = 52; }) (Foo { x = 53; y = 54; }) (Foo { x = 55; y = 56; }) (Foo { x = 57; y = 58; }), Bar { v = vec True True True; w = (True, 0xAABB); z = Foo { x = 3; y = 4; } }); d = (); e = nil; }
      when i == 5 ==> $finish
