Bit#(16) x = 0;
Bit#(8) y = zeroExtend(x);
