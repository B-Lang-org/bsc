module sysParserUninit();
   rule r;
      Bit#(4) x;
      $display(x);
   endrule
endmodule
