function Bit#(t1) f(Bit#(t2) x);
   return zeroExtend(x);
endfunction

