(* synthesize *)
module sysStringTail_Empty();
   rule r;
      $display(stringTail(""));
   endrule
endmodule
