(* synthesize, options="-aggressive-conditions arg" *)
module sysOptionsAttrBad3 ();
endmodule

