module test();

  (* split *)
  rule test;
    $finish(0);
  endrule

endmodule
