package Expr_FieldUpd () where

struct S =
  f :: Bool

x :: S
x = _ { f = True }

