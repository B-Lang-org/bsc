"foo bar \z glurph"
