// Test that an empty list is not ok

(* synthesize *)
(* gate_input_clocks="" *)
module sysGateInputClocks3 (Clock c1, Clock c2, Clock c3) ();
endmodule
