Bit#(5) x;
x = 5 'd 3;
