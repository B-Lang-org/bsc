import TypeclassDupSuperAbstract_Leaf::*;

// Re-export the typeclass, abstractly
export C;

