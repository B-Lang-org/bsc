
interface Ifc;
  (* enable = "" *)
  method Action start(Bool a, Bool b);
endinterface

