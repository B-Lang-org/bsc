package ClassDefResGivenNum () where

class (Foo :: * -> #) a where
    x :: Bool

