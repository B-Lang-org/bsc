-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EUnifyKind.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the EUnifyKind error of the bluespec
-- compiler 
--
-----------------------------------------------------------------------



package EUnifyKind(absval) where

-- import Int

interface Absval  =
         start :: Int a -> Int a 


mkAbsval :: Module (Absval a)
        
mkAbsval = 
        module
           interface
              start x = if x > 0 then
                           x
                        else 
                           negate x  

absval :: Module (Absval 5)
absval = mkAbsval 
