module mkEmptyModuleInterface();
endmodule: mkEmptyModuleInterface
