Bit#(8) x; 
x = 8'b0;