Integer x = 'x;
