(* synthesize *)
module sysPrintType4();

  messageM(printType(typeOf(0)));

endmodule

