package DummyInDefOp () where

(+):: Bool -> Bool -> Bit 12
_ + x = _
