function Action status (Bool a);
action
  while (True)
    $display ("True");
endaction
endfunction : status
