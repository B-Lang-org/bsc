package Zaz;

import XReg::*;

typedef XReg#(a, Bit#(32)) CXReg#(type a);

endpackage
