(* synthesize *)
module sysVerilogElab(Reg#(Bool));
   Reg#(Bool) rg <- mkRegU;
   return rg;
endmodule

