function Bit#(TAdd#(n)) fn(Bit#(n) v1, Bit#(m) v2);
   return {v1, v2};
endfunction
