package StringLit() where

foo :: String
foo = "foo\n"

