function Bool f(Bool something);
  Bool x;
  if (something)
    x = True;
  else
    x = False;
  f = True;
endfunction
