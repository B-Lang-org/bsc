interface Ifc;
  method Action oldname();
endinterface

