
import Foo :: * ;
