export foo;

function a foo(a x) provisos (Bits#(a, sza));
    return (\∘ (unpack, pack))(x);
endfunction: foo

