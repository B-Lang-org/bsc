-- Counter with start value, and upper and lower limits
-- possible to increment and decrement

package Counter (mkCounter, Counter(..)) where

interface Counter a =

   get :: a
   set :: a -> Action

   inc_dec :: Bool -> Action  -- increment if True, otherwise decrement


mkCounter :: (Bits a b, Eq a, Literal a, Arith a) =>
	     a -> a -> a -> Module (Counter a)
mkCounter lower start upper  =
  module

    value_reg :: Reg a <- mkReg start

    interface

      get = value_reg

      set a =
	value_reg := a

      inc_dec up =
	value_reg := if up && value_reg /= upper then
			value_reg + 1
                     else if not up && value_reg /= lower then
                        value_reg - 1
                     else
		        value_reg
