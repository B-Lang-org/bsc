import ReExportItems_Q::*;

// test that the type made it
AB b2 = B;

// test that the variable didn't make it
Bool bOK = b == b2;


