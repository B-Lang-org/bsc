package PolyData(Id(..)) where

data Id = MyId (a -> a)


