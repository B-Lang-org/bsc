(* synthesize *)
module sysEmptyModule ();
endmodule

