(* synthesize, options="aggressive-conditions" *)
module sysOptionsAttrBad1 ();
endmodule

