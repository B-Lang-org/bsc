module ASSIGN1(IN, OUT);
   output OUT;
   input IN;
   assign OUT = IN;
endmodule
