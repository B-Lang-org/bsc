package PolyData2(Id(..)) where

data Id = MyId (a -> a) Integer



