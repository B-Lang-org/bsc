package CDefl () where

import List

x :: Bit a
x = let y :: List a
	y = Nil
    in  fromInteger (length y)

