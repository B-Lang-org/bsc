
// User made a mistake in the syntax
`ifndef (verbosity >= 2)
Bool x = True;
`endif

