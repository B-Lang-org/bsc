
(* synthesize=1, synthesize=0 *)
module sysMultipleAttribModule();
endmodule

