-----------------------------------------------------------------------
-- Project: Bluespec

-- File: ERuleAssertion.bs

-- Author : Amit Grover      <amit@noida.interrasystems.com>

-- Description: This testcase triggers the ERuleAssertion error of the bluespec
-- compiler ("Assertion" failed for rule "RULE")
--
-- Error generated when verilog requested for mkGCD
-----------------------------------------------------------------------



package ERuleAssertion () where

-- import Int

interface GCD =
    start  :: Int 32 -> Int 32 -> Action
    result :: Int 32



mkGCD :: Module GCD
mkGCD =
    module
	x :: Reg (Int 32)
	x <- mkRegU

	y :: Reg (Int 32)
	y <- mkReg 0

        rules
          {-# ASSERT fire when enabled #-}
	  "Swap":
	    when x >= y, y /= 0
	      ==> action
		      x := y
	   	      y := x
          {-# ASSERT fire when enabled #-}
	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0


