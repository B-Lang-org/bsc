package S1;

interface S1#(type aA);
  method aA result(aA c);
  method ActionValue#(aA) check(aA d);
endinterface

endpackage

