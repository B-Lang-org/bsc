module sysAmbigTCon_TAdd (Reg#(Bit#(TAdd#(x,y))));
endmodule
