
Bit#(11) x = 11'h7FF;

Bit#(11) y = -11'h400;

