package DollarColonEqualsPrecedencePretty2 where

foo :: Action -> Action
foo = id

bar :: Reg Bool -> Action
bar r = foo $ (r := False)

