/*
 * comment
 * � with � a � non-ASCII
 * � symbol
 */

export foo;

function a foo(a x);
    return x;
endfunction: foo

