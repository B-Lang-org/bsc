import Vector::*;

Vector#(int, int) initialCoefs;
initialCoefs[0] = 1;
initialCoefs[1] = 1;
initialCoefs[2] = 1;
initialCoefs[3] = 1;
