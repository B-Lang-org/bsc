function Action f();
  action
    f = ?;
  endaction
endfunction
