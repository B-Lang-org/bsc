function Bit#(k) fn (Bit#(m) x, Bit#(n) y)
   provisos (Add#(m, n, Bit#(k)));

   return ?;
endfunction

