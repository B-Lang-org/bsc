// Bug 1336

import "BVI"
   module mkImportModIfc_TooFewArgs(Reg);
      default_clock no_clock;
      default_reset no_reset;
   endmodule

