module sysModDef_PortArg(Bool _, Empty ifc);
  Reg#(Bool) rg <- mkReg(_);
endmodule
