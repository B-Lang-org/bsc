(* synthesize *)
module mkWrongMod ();
endmodule

