package Bug417;
import Bug417::*;
endpackage: Bug417
