interface INonOptionalMethodTypes;
    method m(x, y);
endinterface
