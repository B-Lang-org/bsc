function Bool listy();
  Bool xsss[2][3][5];
  xsss[1][2][3] = True;
  listy = xsss[0][2][4];
endfunction
