import ExportSomeExport::*;

Bool quux;
quux = foo || bar;
