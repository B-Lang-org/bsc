package DegreePrimeVar3(a°) where

a° :: a -> a
a° = id
