package TypeAliasParamGivenNonNumUsedNum () where

type (Foo :: * -> *) a = Bit a

