package ReExportSame_P;

export T(..);

typedef struct {
  Bool f1;
  Bool f2;
 } T;

endpackage
