function Bool f(Bool a);
  Bool x, y;
  x = a;
  return x;
endfunction
