function bit[3:0] f();
  x = 3;
  f = x;
endfunction
