
(* always_ready, always_enabled *)
interface Ifc2;

   (* prefix = "" *)
   method Action m((* port = "VAL" *) Bit#(8) value);
 
endinterface

