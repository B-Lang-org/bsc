`define is 5
`define fs 5
`define full sysFromReal_5_5

`include "FromReal.bsv"
