
(*synthesize*)
module sysInoutProps_UnusedArg #(Inout#(Bit#(32)) io_arg) ();
endmodule

