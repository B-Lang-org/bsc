module mkFoo();
  Bool x = True;
endmodule

