import Vector::*;

(* synthesize *)
module sysRenameResetFail ( (* port="B" *)Vector#(2,Reset) rsts, Empty ifc);
endmodule

