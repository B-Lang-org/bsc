
interface Ifc;
 (* result = "res  ult" *)
 method Bool check ();
endinterface

