module mkFoo();
  rule bogus;
    id(noAction);
  endrule
endmodule
