(* synthesize *)
module mkAbstractDerivePosition();
   primError(?,"should not see");
endmodule
