package TwoArgMissingTwo () where

data Foo a b = Bar a b

x :: Foo
x = _

