package StructDefParamGivenNumUsedNonNum () where

data (Foo :: * -> *) a = Bar a

struct (Baz :: # -> *) b =
    glurph :: Foo b

