package FieldSelectionWithDigit where

x :: Integer
x = foo.bar.0.baz
