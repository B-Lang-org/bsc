import ReExportTestDataConFull::*;

U#(Bool) u = tagged Tag { b1: True, b2: False };
