package ExportAllExportBad() where

foo :: Bool
foo = True

bar :: Bool
bar = False
