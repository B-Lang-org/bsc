package TypeAliasParamGivenTooMany_FromNone () where

type (Foo :: * -> *) = Bit 8

