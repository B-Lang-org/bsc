export はと;

// hiragana are not unicode uppercase letters, so fine for variables

function a はと(a x);
    return id(x);
endfunction: はと

