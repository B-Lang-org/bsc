package TooManyBlockersEsposito(sysTooManyBlockersEsposito) where

-- `Victim' rules are independent and could fire simultaneously
-- were it not for rule `Blocker.'
-- Unlike in the direct test which resorts to using a pri[pars] scheduler,
-- here an Esposito scheduler is produced.  And it allows the victims to
-- fire whenever Blocker is not enabled.

import RegFile
import Vector

type N = 16

sysTooManyBlockersEsposito :: Module Empty
sysTooManyBlockersEsposito =
    module
        arrs :: Vector N (RegFile Bool Bool)
        arrs <- mapM (\_ -> mkRegFileFull) genList
        addRules $ blocker arrs <+> joinRules (map victim arrs)

blocker :: Vector N (RegFile Bool Bool) -> Rules
blocker arrs = rules "Blocker": when True ==> joinActions $ map (\a -> a.upd True True) arrs

victim :: RegFile Bool Bool -> Rules
victim arr = rules "Victim": when True ==> arr.upd True False
