package UTF8BadCons1(鳥(..)) where

-- kanji are not unicode uppercase letters

data 鳥 = 鶴 | 梟

