ActionValue#(Bool) av;
av =
  actionvalue
    return True;
  endactionvalue;
