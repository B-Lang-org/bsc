module mkFoo();
  module mkBar();
  endmodule
endmodule
