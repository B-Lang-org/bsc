package Bug85(mkInterface) where 

import FIFO 

mkInterface :: Bool -> FIFO (Bit 8)
mkInterface b = interface FIFO
		  enq x = noAction
		  first = 12 when b
                  clear = noAction 
                  deq = noAction when b
 
