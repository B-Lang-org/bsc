package StructPat_BadQualField where

import FloatingPoint

fn :: FloatingPoint.Half -> Bit 5
fn (FloatingPoint.Half { sign = True; Foo.exp = e }) = e
fn _ = 0
