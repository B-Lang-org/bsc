
package Foo () where

