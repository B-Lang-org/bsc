Bool data = False;
Bool foreign = False;
Bool in = False;
Bool infix = False;
Bool infixl = False;
Bool infixr = False;
Bool of = False;
Bool prefix = False;
Bool qualified = False;
Bool signature = False;
Bool then = False;
Bool verilog = False;
Bool synthesize = False;
Bool when = False;
Bool where = False;
