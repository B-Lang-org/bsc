package EmptyAction_Layout where

a :: Action
a = action

x :: Integer
x = 17
