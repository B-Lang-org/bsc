typedef union tagged {
   Bool First;
   void Second;
} TaggedUnionSimple;

