(* synthesize, options="-foo" *)
module sysOptionsAttrBad2 ();
endmodule

