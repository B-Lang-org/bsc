module mkFoo();
  rule bogus;
    Bool x;
    x = True;
  endrule
endmodule

