function Bool f();
  Bool x;
  x =True;
  return False;
endfunction
