// Comment

`line(/file/path)

// Comment
