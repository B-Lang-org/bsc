
export Foo::*;

