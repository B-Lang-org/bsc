export 鳩;

// kanji are not unicode uppercase letters, so fine for variables

function a 鳩(a x);
    return id(x);
endfunction: 鳩

