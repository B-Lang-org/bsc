(* synthesize *)
module sysPropDeduce_SubmodUseUnused ();
   Reg#(Bool) r <- mkReg(True);
endmodule

