package Input;

typedef struct {Bit#(129) a;
                Bit#(129) b;
                Bit#(129) bOr;
                Bit#(128) bOr_127;
                Bit#(127) bOr_126;
                Bit#(97) bOr_96;
                Bit#(96) bOr_95;
                Bit#(95) bOr_94;
                Bit#(65) bOr_64;
                Bit#(64) bOr_63;
                Bit#(63) bOr_62;
                Bit#(33) bOr_32;
                Bit#(32) bOr_31;
                Bit#(31) bOr_30;
                Bit#(2) bOr_1;
                Bit#(1) bOr_0;
                Bit#(129) bAnd;
                Bit#(128) bAnd_127;
                Bit#(127) bAnd_126;
                Bit#(97) bAnd_96;
                Bit#(96) bAnd_95;
                Bit#(95) bAnd_94;
                Bit#(65) bAnd_64;
                Bit#(64) bAnd_63;
                Bit#(63) bAnd_62;
                Bit#(33) bAnd_32;
                Bit#(32) bAnd_31;
                Bit#(31) bAnd_30;
                Bit#(2) bAnd_1;
                Bit#(1) bAnd_0;
                Bit#(129) bInv;
                Bit#(128) bInv_127;
                Bit#(127) bInv_126;
                Bit#(97) bInv_96;
                Bit#(96) bInv_95;
                Bit#(95) bInv_94;
                Bit#(65) bInv_64;
                Bit#(64) bInv_63;
                Bit#(63) bInv_62;
                Bit#(33) bInv_32;
                Bit#(32) bInv_31;
                Bit#(31) bInv_30;
                Bit#(2) bInv_1;
                Bit#(1) bInv_0;
                Bit#(129) bXor;
                Bit#(128) bXor_127;
                Bit#(127) bXor_126;
                Bit#(97) bXor_96;
                Bit#(96) bXor_95;
                Bit#(95) bXor_94;
                Bit#(65) bXor_64;
                Bit#(64) bXor_63;
                Bit#(63) bXor_62;
                Bit#(33) bXor_32;
                Bit#(32) bXor_31;
                Bit#(31) bXor_30;
                Bit#(2) bXor_1;
                Bit#(1) bXor_0;
                Bit#(129) bXnor;
                Bit#(128) bXnor_127;
                Bit#(127) bXnor_126;
                Bit#(97) bXnor_96;
                Bit#(96) bXnor_95;
                Bit#(95) bXnor_94;
                Bit#(65) bXnor_64;
                Bit#(64) bXnor_63;
                Bit#(63) bXnor_62;
                Bit#(33) bXnor_32;
                Bit#(32) bXnor_31;
                Bit#(31) bXnor_30;
                Bit#(2) bXnor_1;
                Bit#(1) bXnor_0;
				} Inputs deriving(Bits,Eq);

endpackage : Input 
