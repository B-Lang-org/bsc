package StructDefResGivenNum () where

struct (Foo :: #) =
    x :: Bool

