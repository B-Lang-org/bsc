import Prelude :: *;
