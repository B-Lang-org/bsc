package TypeAliasParamGivenTooFew () where

type (Foo :: * -> *) a b = Tuple2 a b

