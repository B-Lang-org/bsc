package TypeAliasPartialAppWithConflictingKindSig () where

type (Foo :: * -> *) = Bit

