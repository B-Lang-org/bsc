module mkEmptyRule(Empty);
    rule emptyrule;
    endrule
endmodule: mkEmptyRule
