package RecDeriveDataOneArg () where

data Foo = F Foo deriving (Eq)

