module mkFoo();
  Reg#(Bool) r();
  mkReg#(True) the_r(r);
endmodule
