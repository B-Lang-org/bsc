package FFReadTest(sysFFReadTest) where

sysFFReadTest :: Module Empty
sysFFReadTest = 
  module
    r :: Reg (Bit 16) <- mkReg 7
    done :: Reg (Bool) <- mkReg False

    rules 
      when done ==> $finish 0
      when not done ==> 
        action
          displayHex r
          done := True