package Displayable(Displayable(..)) where

class Displayable a where
   display :: a -> Action

instance (Bits a sa) => Displayable a
   where
     display a = $display "Bits %h" a
