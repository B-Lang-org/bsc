// Comment

`line(/file/path,4,1,0
