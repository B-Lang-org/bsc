package StructDefFieldIsNum () where

struct Foo =
    bar :: 12

