
interface Ifc;
 method Action check ((* port="arg" *) (* port="arg" *)Bool x);
endinterface

