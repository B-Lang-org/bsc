import TypeclassDup_Leaf::*;

export Expose(..);

