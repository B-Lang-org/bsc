(* synthesize *)
module sysInvalid_Bit_Bin ();
   Reg#(Bit#(4)) rg <- mkReg('b10101);
endmodule
