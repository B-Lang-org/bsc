// This is the original example for Bug 991.

typedef union tagged {
   a T1;
} U#(numeric type a);

