Integer test = True;

(* synthesize *)
module sysDefErrorRecovery();

  rule test;
    $display("Test passed\n");
  endrule

endmodule
