-----------------------------------------------------------------------
-- Project: Bluespec

-- File: EUnify1.bs

-- Author : Nitin Chand Rahul      <ncr@noida.interrasystems.com>

-- Description: This testcase triggers a Type error (EUnify)

-- Error Message : bsc EUnify1.bs
-- bsc: Compilation errors:
-- "EUnify1.bs", line 54, column 12, Type error at:
-- start

-- Expected type:
-- Prelude.Action

-- Inferred type:
-- Int.Int 32 -> Int.Int 32 -> Prelude.Action
-----------------------------------------------------------------------

package EUnify1 (EUnify1(..), mkEUnify1) where

-- import Int

interface EUnify1 =
    start  :: Action
    result :: Int 32


mkEUnify1 :: Module EUnify1
mkEUnify1 =
    module

        x :: Reg (Int 32)
        x <- mkReg 0

	y :: Reg (Int 32)
	y <- mkReg 0
       
        rules
	  "Swap":
	    when x > y, y /= 0
	      ==> action
		      x := y
		      y := x

	  "Subtract":
	    when x <= y, y /= 0
	      ==> action
		      y := y - x

        interface
	    start ix iy = action
	                      x := ix
	                      y := iy
	                  when y == 0
	    result = x when y == 0
