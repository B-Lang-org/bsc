package Primitive () where

primitive _ :: Bit 1

