function Bool f(a#(n) y);
  a x = ?;
  return True;
endfunction


