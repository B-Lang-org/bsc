package Design_seq ;

interface Design_seq_IFC #(parameter type a,parameter type b);
    method Action seq(a namea ,a nameb);
    method b speed();
endinterface:  Design_seq_IFC

endpackage: Design_seq

